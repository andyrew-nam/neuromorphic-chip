`timescale 1ns / 1ps

module hazard_detector_nn (
    input wire clk,
    input wire rst,
    input wire start,
    input wire [7:0] image_pixels [0:207],  // 208 pixels, 8-bit grayscale
    output reg done,
    output reg [15:0] outputs [0:14]        // 15 outputs Q8.8 fixed-point
);

    // Sizes
    localparam IN_SIZE = 208;
    localparam H1_SIZE = 128;
    localparam H2_SIZE = 64;
    localparam OUT_SIZE = 15;

    // Fixed-point Q8.8 signed format
    // 16 bits: [15] sign, [14:8] integer, [7:0] fraction

    // State machine states
    typedef enum reg [3:0] {  // Changed to 4 bits to accommodate new state
        IDLE,
        LAYER1_NEURON,
        LAYER1_MAC,
        LAYER1_RELU,
        LAYER2_NEURON,
        LAYER2_MAC,
        LAYER2_RELU,
        LAYER3_NEURON,
        LAYER3_MAC,
        LAYER3_SIGMOID,
        COPY_OUTPUTS,  // New state for copying outputs
        DONE_STATE
    } state_t;

    state_t state;

    // Counters for neurons and inputs
    reg [7:0] neuron_idx;    // Enough for max 128 neurons
    reg [7:0] input_idx;

    // Accumulator for MAC (32-bit signed to avoid overflow)
    reg signed [31:0] acc;

    // Intermediate neuron output storage
    reg signed [15:0] layer1_out [0:H1_SIZE-1];
    reg signed [15:0] layer2_out [0:H2_SIZE-1];

    // Weights and biases
    reg signed [15:0] fc1_weights [0:H1_SIZE-1][0:IN_SIZE-1];
    reg signed [15:0] fc1_biases  [0:H1_SIZE-1];

    reg signed [15:0] fc2_weights [0:H2_SIZE-1][0:H1_SIZE-1];
    reg signed [15:0] fc2_biases  [0:H2_SIZE-1];

    reg signed [15:0] fc3_weights [0:OUT_SIZE-1][0:H2_SIZE-1];
    reg signed [15:0] fc3_biases  [0:OUT_SIZE-1];

    // Output registers
    reg signed [15:0] fc3_out [0:OUT_SIZE-1];

    // ReLU activation
    function signed [15:0] relu;
        input signed [31:0] x;
        begin
            if (x < 0)
                relu = 0;
            else if (x > 32767)
                relu = 32767;
            else
                relu = x[15:0]; // Keep lower 16 bits after MAC shift (you may need shift)
        end
    endfunction

    // Sigmoid approximation (hard sigmoid)
    function signed [15:0] sigmoid_approx;
        input signed [15:0] x;
        reg signed [15:0] val;
        begin
            // scale input from Q8.8 to approx range and clip
            // simple: f(x) = max(0, min(1, 0.5 + x/4))
            val = 16'd128 + (x >>> 2);
            if (val < 0)
                sigmoid_approx = 0;
            else if (val > 16'd256)
                sigmoid_approx = 16'd256;
            else
                sigmoid_approx = val;
        end
    endfunction

    // Main sequential logic
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            done <= 0;
            neuron_idx <= 0;
            input_idx <= 0;
            acc <= 0;
        end else begin
            case (state)

                IDLE: begin
                    done <= 0;
                    neuron_idx <= 0;
                    input_idx <= 0;
                    acc <= 0;
                    if (start)
                        state <= LAYER1_NEURON;
                end

                // Layer 1: compute each neuron MAC sequentially
                LAYER1_NEURON: begin
                    acc <= (fc1_biases[neuron_idx] <<< 8);  // bias scaled to Q16.16 for accumulation
                    input_idx <= 0;
                    state <= LAYER1_MAC;
                end

                LAYER1_MAC: begin
                    acc <= acc + $signed(fc1_weights[neuron_idx][input_idx]) * $signed({8'd0, image_pixels[input_idx]});
                    if (input_idx == IN_SIZE - 1)
                        state <= LAYER1_RELU;
                    else
                        input_idx <= input_idx + 1;
                end

                LAYER1_RELU: begin
                    layer1_out[neuron_idx] <= relu(acc >>> 8); // shift back from Q16.16 to Q8.8
                    if (neuron_idx == H1_SIZE - 1) begin
                        neuron_idx <= 0;
                        state <= LAYER2_NEURON;
                    end else
                        neuron_idx <= neuron_idx + 1;
                end

                // Layer 2: same sequential MAC for hidden layer 2
                LAYER2_NEURON: begin
                    acc <= (fc2_biases[neuron_idx] <<< 8);
                    input_idx <= 0;
                    state <= LAYER2_MAC;
                end

                LAYER2_MAC: begin
                    acc <= acc + $signed(fc2_weights[neuron_idx][input_idx]) * $signed(layer1_out[input_idx]);
                    if (input_idx == H1_SIZE - 1)
                        state <= LAYER2_RELU;
                    else
                        input_idx <= input_idx + 1;
                end

                LAYER2_RELU: begin
                    layer2_out[neuron_idx] <= relu(acc >>> 8);
                    if (neuron_idx == H2_SIZE - 1) begin
                        neuron_idx <= 0;
                        state <= LAYER3_NEURON;
                    end else
                        neuron_idx <= neuron_idx + 1;
                end

                // Layer 3: output layer neurons
                LAYER3_NEURON: begin
                    acc <= (fc3_biases[neuron_idx] <<< 8);
                    input_idx <= 0;
                    state <= LAYER3_MAC;
                end

                LAYER3_MAC: begin
                    acc <= acc + $signed(fc3_weights[neuron_idx][input_idx]) * $signed(layer2_out[input_idx]);
                    if (input_idx == H2_SIZE - 1)
                        state <= LAYER3_SIGMOID;
                    else
                        input_idx <= input_idx + 1;
                end

                LAYER3_SIGMOID: begin
                    fc3_out[neuron_idx] <= sigmoid_approx(acc[23:8]); // use middle bits for Q8.8
                    if (neuron_idx == OUT_SIZE - 1) begin
                        neuron_idx <= 0;  // Reset counter for copying outputs
                        state <= COPY_OUTPUTS;
                    end else
                        neuron_idx <= neuron_idx + 1;
                end

                // New state to copy outputs sequentially
                COPY_OUTPUTS: begin
                    outputs[neuron_idx] <= fc3_out[neuron_idx];
                    if (neuron_idx == OUT_SIZE - 1) begin
                        done <= 1;
                        state <= DONE_STATE;
                    end else
                        neuron_idx <= neuron_idx + 1;
                end

                DONE_STATE: begin
                    if (!start)
                        state <= IDLE;
                end

                default: state <= IDLE;
            endcase
        end
    end

    initial begin
        // Auto-generated Verilog weight initialization (Q8.8 fixed-point, 16-bit signed)
        // Copy these lines into your Verilog module's initial block
        
        // fc1 weights
        fc1_weights[0][0] = 16'sd8;
        fc1_weights[0][1] = 16'sd-6;
        fc1_weights[0][2] = 16'sd-12;
        fc1_weights[0][3] = 16'sd-11;
        fc1_weights[0][4] = 16'sd-48;
        fc1_weights[0][5] = 16'sd-20;
        fc1_weights[0][6] = 16'sd-10;
        fc1_weights[0][7] = 16'sd-54;
        fc1_weights[0][8] = 16'sd-5;
        fc1_weights[0][9] = 16'sd-2;
        fc1_weights[0][10] = 16'sd-18;
        fc1_weights[0][11] = 16'sd-41;
        fc1_weights[0][12] = 16'sd48;
        fc1_weights[0][13] = 16'sd32;
        fc1_weights[0][14] = 16'sd-22;
        fc1_weights[0][15] = 16'sd-39;
        fc1_weights[0][16] = 16'sd-4;
        fc1_weights[0][17] = 16'sd70;
        fc1_weights[0][18] = 16'sd49;
        fc1_weights[0][19] = 16'sd19;
        fc1_weights[0][20] = 16'sd-30;
        fc1_weights[0][21] = 16'sd-49;
        fc1_weights[0][22] = 16'sd-26;
        fc1_weights[0][23] = 16'sd31;
        fc1_weights[0][24] = 16'sd-44;
        fc1_weights[0][25] = 16'sd4;
        fc1_weights[0][26] = 16'sd42;
        fc1_weights[0][27] = 16'sd-6;
        fc1_weights[0][28] = 16'sd7;
        fc1_weights[0][29] = 16'sd16;
        fc1_weights[0][30] = 16'sd-5;
        fc1_weights[0][31] = 16'sd1;
        fc1_weights[0][32] = 16'sd9;
        fc1_weights[0][33] = 16'sd5;
        fc1_weights[0][34] = 16'sd-7;
        fc1_weights[0][35] = 16'sd-13;
        fc1_weights[0][36] = 16'sd-66;
        fc1_weights[0][37] = 16'sd-49;
        fc1_weights[0][38] = 16'sd-7;
        fc1_weights[0][39] = 16'sd-17;
        fc1_weights[0][40] = 16'sd-87;
        fc1_weights[0][41] = 16'sd-7;
        fc1_weights[0][42] = 16'sd55;
        fc1_weights[0][43] = 16'sd37;
        fc1_weights[0][44] = 16'sd17;
        fc1_weights[0][45] = 16'sd-10;
        fc1_weights[0][46] = 16'sd61;
        fc1_weights[0][47] = 16'sd3;
        fc1_weights[0][48] = 16'sd-18;
        fc1_weights[0][49] = 16'sd6;
        fc1_weights[0][50] = 16'sd34;
        fc1_weights[0][51] = 16'sd57;
        fc1_weights[0][52] = 16'sd53;
        fc1_weights[0][53] = 16'sd7;
        fc1_weights[0][54] = 16'sd-8;
        fc1_weights[0][55] = 16'sd54;
        fc1_weights[0][56] = 16'sd7;
        fc1_weights[0][57] = 16'sd0;
        fc1_weights[0][58] = 16'sd-21;
        fc1_weights[0][59] = 16'sd-52;
        fc1_weights[0][60] = 16'sd-25;
        fc1_weights[0][61] = 16'sd13;
        fc1_weights[0][62] = 16'sd-62;
        fc1_weights[0][63] = 16'sd-58;
        fc1_weights[0][64] = 16'sd-88;
        fc1_weights[0][65] = 16'sd-45;
        fc1_weights[0][66] = 16'sd-49;
        fc1_weights[0][67] = 16'sd15;
        fc1_weights[0][68] = 16'sd-24;
        fc1_weights[0][69] = 16'sd58;
        fc1_weights[0][70] = 16'sd13;
        fc1_weights[0][71] = 16'sd38;
        fc1_weights[0][72] = 16'sd-8;
        fc1_weights[0][73] = 16'sd55;
        fc1_weights[0][74] = 16'sd16;
        fc1_weights[0][75] = 16'sd6;
        fc1_weights[0][76] = 16'sd-17;
        fc1_weights[0][77] = 16'sd7;
        fc1_weights[0][78] = 16'sd38;
        fc1_weights[0][79] = 16'sd-25;
        fc1_weights[0][80] = 16'sd18;
        fc1_weights[0][81] = 16'sd46;
        fc1_weights[0][82] = 16'sd-23;
        fc1_weights[0][83] = 16'sd36;
        fc1_weights[0][84] = 16'sd30;
        fc1_weights[0][85] = 16'sd6;
        fc1_weights[0][86] = 16'sd22;
        fc1_weights[0][87] = 16'sd17;
        fc1_weights[0][88] = 16'sd85;
        fc1_weights[0][89] = 16'sd-2;
        fc1_weights[0][90] = 16'sd-69;
        fc1_weights[0][91] = 16'sd-66;
        fc1_weights[0][92] = 16'sd-10;
        fc1_weights[0][93] = 16'sd8;
        fc1_weights[0][94] = 16'sd17;
        fc1_weights[0][95] = 16'sd-25;
        fc1_weights[0][96] = 16'sd-2;
        fc1_weights[0][97] = 16'sd-3;
        fc1_weights[0][98] = 16'sd5;
        fc1_weights[0][99] = 16'sd11;
        fc1_weights[0][100] = 16'sd2;
        fc1_weights[0][101] = 16'sd11;
        fc1_weights[0][102] = 16'sd21;
        fc1_weights[0][103] = 16'sd77;
        fc1_weights[0][104] = 16'sd-7;
        fc1_weights[0][105] = 16'sd22;
        fc1_weights[0][106] = 16'sd27;
        fc1_weights[0][107] = 16'sd49;
        fc1_weights[0][108] = 16'sd2;
        fc1_weights[0][109] = 16'sd22;
        fc1_weights[0][110] = 16'sd-18;
        fc1_weights[0][111] = 16'sd-13;
        fc1_weights[0][112] = 16'sd-1;
        fc1_weights[0][113] = 16'sd52;
        fc1_weights[0][114] = 16'sd21;
        fc1_weights[0][115] = 16'sd-4;
        fc1_weights[0][116] = 16'sd22;
        fc1_weights[0][117] = 16'sd-17;
        fc1_weights[0][118] = 16'sd-18;
        fc1_weights[0][119] = 16'sd30;
        fc1_weights[0][120] = 16'sd50;
        fc1_weights[0][121] = 16'sd-9;
        fc1_weights[0][122] = 16'sd-15;
        fc1_weights[0][123] = 16'sd55;
        fc1_weights[0][124] = 16'sd53;
        fc1_weights[0][125] = 16'sd57;
        fc1_weights[0][126] = 16'sd108;
        fc1_weights[0][127] = 16'sd27;
        fc1_weights[0][128] = 16'sd32;
        fc1_weights[0][129] = 16'sd160;
        fc1_weights[0][130] = 16'sd-18;
        fc1_weights[0][131] = 16'sd-34;
        fc1_weights[0][132] = 16'sd24;
        fc1_weights[0][133] = 16'sd1;
        fc1_weights[0][134] = 16'sd-41;
        fc1_weights[0][135] = 16'sd-26;
        fc1_weights[0][136] = 16'sd12;
        fc1_weights[0][137] = 16'sd-71;
        fc1_weights[0][138] = 16'sd-121;
        fc1_weights[0][139] = 16'sd-84;
        fc1_weights[0][140] = 16'sd0;
        fc1_weights[0][141] = 16'sd-42;
        fc1_weights[0][142] = 16'sd-15;
        fc1_weights[0][143] = 16'sd34;
        fc1_weights[0][144] = 16'sd13;
        fc1_weights[0][145] = 16'sd14;
        fc1_weights[0][146] = 16'sd15;
        fc1_weights[0][147] = 16'sd30;
        fc1_weights[0][148] = 16'sd46;
        fc1_weights[0][149] = 16'sd37;
        fc1_weights[0][150] = 16'sd49;
        fc1_weights[0][151] = 16'sd37;
        fc1_weights[0][152] = 16'sd16;
        fc1_weights[0][153] = 16'sd5;
        fc1_weights[0][154] = 16'sd2;
        fc1_weights[0][155] = 16'sd29;
        fc1_weights[0][156] = 16'sd60;
        fc1_weights[0][157] = 16'sd24;
        fc1_weights[0][158] = 16'sd44;
        fc1_weights[0][159] = 16'sd12;
        fc1_weights[0][160] = 16'sd-23;
        fc1_weights[0][161] = 16'sd-19;
        fc1_weights[0][162] = 16'sd-68;
        fc1_weights[0][163] = 16'sd38;
        fc1_weights[0][164] = 16'sd20;
        fc1_weights[0][165] = 16'sd17;
        fc1_weights[0][166] = 16'sd-33;
        fc1_weights[0][167] = 16'sd-43;
        fc1_weights[0][168] = 16'sd-28;
        fc1_weights[0][169] = 16'sd6;
        fc1_weights[0][170] = 16'sd-27;
        fc1_weights[0][171] = 16'sd-92;
        fc1_weights[0][172] = 16'sd-52;
        fc1_weights[0][173] = 16'sd-48;
        fc1_weights[0][174] = 16'sd-32;
        fc1_weights[0][175] = 16'sd17;
        fc1_weights[0][176] = 16'sd21;
        fc1_weights[0][177] = 16'sd-12;
        fc1_weights[0][178] = 16'sd60;
        fc1_weights[0][179] = 16'sd11;
        fc1_weights[0][180] = 16'sd77;
        fc1_weights[0][181] = 16'sd15;
        fc1_weights[0][182] = 16'sd-45;
        fc1_weights[0][183] = 16'sd-18;
        fc1_weights[0][184] = 16'sd0;
        fc1_weights[0][185] = 16'sd-62;
        fc1_weights[0][186] = 16'sd-43;
        fc1_weights[0][187] = 16'sd-12;
        fc1_weights[0][188] = 16'sd-25;
        fc1_weights[0][189] = 16'sd32;
        fc1_weights[0][190] = 16'sd40;
        fc1_weights[0][191] = 16'sd-27;
        fc1_weights[0][192] = 16'sd62;
        fc1_weights[0][193] = 16'sd23;
        fc1_weights[0][194] = 16'sd-2;
        fc1_weights[0][195] = 16'sd5;
        fc1_weights[0][196] = 16'sd42;
        fc1_weights[0][197] = 16'sd-80;
        fc1_weights[0][198] = 16'sd-57;
        fc1_weights[0][199] = 16'sd-35;
        fc1_weights[0][200] = 16'sd-50;
        fc1_weights[0][201] = 16'sd11;
        fc1_weights[0][202] = 16'sd-74;
        fc1_weights[0][203] = 16'sd-38;
        fc1_weights[0][204] = 16'sd-52;
        fc1_weights[0][205] = 16'sd-30;
        fc1_weights[0][206] = 16'sd11;
        fc1_weights[0][207] = 16'sd36;
        fc1_weights[1][0] = 16'sd68;
        fc1_weights[1][1] = 16'sd-38;
        fc1_weights[1][2] = 16'sd16;
        fc1_weights[1][3] = 16'sd52;
        fc1_weights[1][4] = 16'sd49;
        fc1_weights[1][5] = 16'sd13;
        fc1_weights[1][6] = 16'sd48;
        fc1_weights[1][7] = 16'sd-8;
        fc1_weights[1][8] = 16'sd36;
        fc1_weights[1][9] = 16'sd133;
        fc1_weights[1][10] = 16'sd54;
        fc1_weights[1][11] = 16'sd77;
        fc1_weights[1][12] = 16'sd97;
        fc1_weights[1][13] = 16'sd-15;
        fc1_weights[1][14] = 16'sd87;
        fc1_weights[1][15] = 16'sd-17;
        fc1_weights[1][16] = 16'sd-51;
        fc1_weights[1][17] = 16'sd-31;
        fc1_weights[1][18] = 16'sd8;
        fc1_weights[1][19] = 16'sd25;
        fc1_weights[1][20] = 16'sd30;
        fc1_weights[1][21] = 16'sd22;
        fc1_weights[1][22] = 16'sd-2;
        fc1_weights[1][23] = 16'sd2;
        fc1_weights[1][24] = 16'sd24;
        fc1_weights[1][25] = 16'sd-52;
        fc1_weights[1][26] = 16'sd73;
        fc1_weights[1][27] = 16'sd34;
        fc1_weights[1][28] = 16'sd33;
        fc1_weights[1][29] = 16'sd-79;
        fc1_weights[1][30] = 16'sd-59;
        fc1_weights[1][31] = 16'sd-99;
        fc1_weights[1][32] = 16'sd-45;
        fc1_weights[1][33] = 16'sd79;
        fc1_weights[1][34] = 16'sd-31;
        fc1_weights[1][35] = 16'sd42;
        fc1_weights[1][36] = 16'sd-53;
        fc1_weights[1][37] = 16'sd40;
        fc1_weights[1][38] = 16'sd35;
        fc1_weights[1][39] = 16'sd98;
        fc1_weights[1][40] = 16'sd-26;
        fc1_weights[1][41] = 16'sd83;
        fc1_weights[1][42] = 16'sd52;
        fc1_weights[1][43] = 16'sd-8;
        fc1_weights[1][44] = 16'sd53;
        fc1_weights[1][45] = 16'sd45;
        fc1_weights[1][46] = 16'sd27;
        fc1_weights[1][47] = 16'sd-1;
        fc1_weights[1][48] = 16'sd24;
        fc1_weights[1][49] = 16'sd-96;
        fc1_weights[1][50] = 16'sd27;
        fc1_weights[1][51] = 16'sd55;
        fc1_weights[1][52] = 16'sd-2;
        fc1_weights[1][53] = 16'sd-21;
        fc1_weights[1][54] = 16'sd-17;
        fc1_weights[1][55] = 16'sd-4;
        fc1_weights[1][56] = 16'sd43;
        fc1_weights[1][57] = 16'sd47;
        fc1_weights[1][58] = 16'sd11;
        fc1_weights[1][59] = 16'sd33;
        fc1_weights[1][60] = 16'sd-96;
        fc1_weights[1][61] = 16'sd-28;
        fc1_weights[1][62] = 16'sd-15;
        fc1_weights[1][63] = 16'sd-37;
        fc1_weights[1][64] = 16'sd-44;
        fc1_weights[1][65] = 16'sd105;
        fc1_weights[1][66] = 16'sd-88;
        fc1_weights[1][67] = 16'sd90;
        fc1_weights[1][68] = 16'sd43;
        fc1_weights[1][69] = 16'sd-55;
        fc1_weights[1][70] = 16'sd-1;
        fc1_weights[1][71] = 16'sd34;
        fc1_weights[1][72] = 16'sd22;
        fc1_weights[1][73] = 16'sd16;
        fc1_weights[1][74] = 16'sd-17;
        fc1_weights[1][75] = 16'sd-13;
        fc1_weights[1][76] = 16'sd-37;
        fc1_weights[1][77] = 16'sd-3;
        fc1_weights[1][78] = 16'sd45;
        fc1_weights[1][79] = 16'sd-63;
        fc1_weights[1][80] = 16'sd-3;
        fc1_weights[1][81] = 16'sd-3;
        fc1_weights[1][82] = 16'sd5;
        fc1_weights[1][83] = 16'sd10;
        fc1_weights[1][84] = 16'sd-8;
        fc1_weights[1][85] = 16'sd25;
        fc1_weights[1][86] = 16'sd-76;
        fc1_weights[1][87] = 16'sd-17;
        fc1_weights[1][88] = 16'sd-88;
        fc1_weights[1][89] = 16'sd-90;
        fc1_weights[1][90] = 16'sd-44;
        fc1_weights[1][91] = 16'sd-86;
        fc1_weights[1][92] = 16'sd-109;
        fc1_weights[1][93] = 16'sd-17;
        fc1_weights[1][94] = 16'sd-65;
        fc1_weights[1][95] = 16'sd-73;
        fc1_weights[1][96] = 16'sd-11;
        fc1_weights[1][97] = 16'sd-42;
        fc1_weights[1][98] = 16'sd-26;
        fc1_weights[1][99] = 16'sd-8;
        fc1_weights[1][100] = 16'sd-40;
        fc1_weights[1][101] = 16'sd-23;
        fc1_weights[1][102] = 16'sd22;
        fc1_weights[1][103] = 16'sd24;
        fc1_weights[1][104] = 16'sd-3;
        fc1_weights[1][105] = 16'sd23;
        fc1_weights[1][106] = 16'sd-18;
        fc1_weights[1][107] = 16'sd0;
        fc1_weights[1][108] = 16'sd-10;
        fc1_weights[1][109] = 16'sd-8;
        fc1_weights[1][110] = 16'sd-35;
        fc1_weights[1][111] = 16'sd-26;
        fc1_weights[1][112] = 16'sd-74;
        fc1_weights[1][113] = 16'sd-23;
        fc1_weights[1][114] = 16'sd9;
        fc1_weights[1][115] = 16'sd21;
        fc1_weights[1][116] = 16'sd75;
        fc1_weights[1][117] = 16'sd-44;
        fc1_weights[1][118] = 16'sd66;
        fc1_weights[1][119] = 16'sd49;
        fc1_weights[1][120] = 16'sd-23;
        fc1_weights[1][121] = 16'sd-52;
        fc1_weights[1][122] = 16'sd-49;
        fc1_weights[1][123] = 16'sd-53;
        fc1_weights[1][124] = 16'sd-3;
        fc1_weights[1][125] = 16'sd7;
        fc1_weights[1][126] = 16'sd-22;
        fc1_weights[1][127] = 16'sd-38;
        fc1_weights[1][128] = 16'sd10;
        fc1_weights[1][129] = 16'sd45;
        fc1_weights[1][130] = 16'sd-1;
        fc1_weights[1][131] = 16'sd6;
        fc1_weights[1][132] = 16'sd2;
        fc1_weights[1][133] = 16'sd33;
        fc1_weights[1][134] = 16'sd-32;
        fc1_weights[1][135] = 16'sd-12;
        fc1_weights[1][136] = 16'sd33;
        fc1_weights[1][137] = 16'sd27;
        fc1_weights[1][138] = 16'sd-20;
        fc1_weights[1][139] = 16'sd88;
        fc1_weights[1][140] = 16'sd19;
        fc1_weights[1][141] = 16'sd40;
        fc1_weights[1][142] = 16'sd11;
        fc1_weights[1][143] = 16'sd98;
        fc1_weights[1][144] = 16'sd-50;
        fc1_weights[1][145] = 16'sd37;
        fc1_weights[1][146] = 16'sd14;
        fc1_weights[1][147] = 16'sd44;
        fc1_weights[1][148] = 16'sd21;
        fc1_weights[1][149] = 16'sd52;
        fc1_weights[1][150] = 16'sd-2;
        fc1_weights[1][151] = 16'sd4;
        fc1_weights[1][152] = 16'sd19;
        fc1_weights[1][153] = 16'sd-57;
        fc1_weights[1][154] = 16'sd-47;
        fc1_weights[1][155] = 16'sd-30;
        fc1_weights[1][156] = 16'sd-23;
        fc1_weights[1][157] = 16'sd-13;
        fc1_weights[1][158] = 16'sd19;
        fc1_weights[1][159] = 16'sd24;
        fc1_weights[1][160] = 16'sd66;
        fc1_weights[1][161] = 16'sd69;
        fc1_weights[1][162] = 16'sd-33;
        fc1_weights[1][163] = 16'sd12;
        fc1_weights[1][164] = 16'sd45;
        fc1_weights[1][165] = 16'sd59;
        fc1_weights[1][166] = 16'sd36;
        fc1_weights[1][167] = 16'sd54;
        fc1_weights[1][168] = 16'sd2;
        fc1_weights[1][169] = 16'sd58;
        fc1_weights[1][170] = 16'sd39;
        fc1_weights[1][171] = 16'sd77;
        fc1_weights[1][172] = 16'sd-25;
        fc1_weights[1][173] = 16'sd26;
        fc1_weights[1][174] = 16'sd36;
        fc1_weights[1][175] = 16'sd66;
        fc1_weights[1][176] = 16'sd5;
        fc1_weights[1][177] = 16'sd-66;
        fc1_weights[1][178] = 16'sd36;
        fc1_weights[1][179] = 16'sd-15;
        fc1_weights[1][180] = 16'sd-48;
        fc1_weights[1][181] = 16'sd21;
        fc1_weights[1][182] = 16'sd-43;
        fc1_weights[1][183] = 16'sd-41;
        fc1_weights[1][184] = 16'sd-8;
        fc1_weights[1][185] = 16'sd-69;
        fc1_weights[1][186] = 16'sd-26;
        fc1_weights[1][187] = 16'sd-55;
        fc1_weights[1][188] = 16'sd-57;
        fc1_weights[1][189] = 16'sd11;
        fc1_weights[1][190] = 16'sd-11;
        fc1_weights[1][191] = 16'sd-55;
        fc1_weights[1][192] = 16'sd-17;
        fc1_weights[1][193] = 16'sd19;
        fc1_weights[1][194] = 16'sd9;
        fc1_weights[1][195] = 16'sd-22;
        fc1_weights[1][196] = 16'sd39;
        fc1_weights[1][197] = 16'sd14;
        fc1_weights[1][198] = 16'sd94;
        fc1_weights[1][199] = 16'sd-7;
        fc1_weights[1][200] = 16'sd-33;
        fc1_weights[1][201] = 16'sd48;
        fc1_weights[1][202] = 16'sd-77;
        fc1_weights[1][203] = 16'sd-117;
        fc1_weights[1][204] = 16'sd-64;
        fc1_weights[1][205] = 16'sd-24;
        fc1_weights[1][206] = 16'sd-14;
        fc1_weights[1][207] = 16'sd-9;
        fc1_weights[2][0] = 16'sd21;
        fc1_weights[2][1] = 16'sd-38;
        fc1_weights[2][2] = 16'sd-28;
        fc1_weights[2][3] = 16'sd-22;
        fc1_weights[2][4] = 16'sd-14;
        fc1_weights[2][5] = 16'sd31;
        fc1_weights[2][6] = 16'sd8;
        fc1_weights[2][7] = 16'sd18;
        fc1_weights[2][8] = 16'sd-82;
        fc1_weights[2][9] = 16'sd-72;
        fc1_weights[2][10] = 16'sd-51;
        fc1_weights[2][11] = 16'sd-85;
        fc1_weights[2][12] = 16'sd-59;
        fc1_weights[2][13] = 16'sd-5;
        fc1_weights[2][14] = 16'sd99;
        fc1_weights[2][15] = 16'sd82;
        fc1_weights[2][16] = 16'sd64;
        fc1_weights[2][17] = 16'sd41;
        fc1_weights[2][18] = 16'sd71;
        fc1_weights[2][19] = 16'sd-41;
        fc1_weights[2][20] = 16'sd-21;
        fc1_weights[2][21] = 16'sd10;
        fc1_weights[2][22] = 16'sd30;
        fc1_weights[2][23] = 16'sd-41;
        fc1_weights[2][24] = 16'sd37;
        fc1_weights[2][25] = 16'sd28;
        fc1_weights[2][26] = 16'sd30;
        fc1_weights[2][27] = 16'sd-87;
        fc1_weights[2][28] = 16'sd-45;
        fc1_weights[2][29] = 16'sd-14;
        fc1_weights[2][30] = 16'sd12;
        fc1_weights[2][31] = 16'sd10;
        fc1_weights[2][32] = 16'sd12;
        fc1_weights[2][33] = 16'sd-32;
        fc1_weights[2][34] = 16'sd-61;
        fc1_weights[2][35] = 16'sd-43;
        fc1_weights[2][36] = 16'sd-27;
        fc1_weights[2][37] = 16'sd-22;
        fc1_weights[2][38] = 16'sd-26;
        fc1_weights[2][39] = 16'sd-41;
        fc1_weights[2][40] = 16'sd139;
        fc1_weights[2][41] = 16'sd104;
        fc1_weights[2][42] = 16'sd5;
        fc1_weights[2][43] = 16'sd81;
        fc1_weights[2][44] = 16'sd47;
        fc1_weights[2][45] = 16'sd-10;
        fc1_weights[2][46] = 16'sd33;
        fc1_weights[2][47] = 16'sd-62;
        fc1_weights[2][48] = 16'sd21;
        fc1_weights[2][49] = 16'sd31;
        fc1_weights[2][50] = 16'sd39;
        fc1_weights[2][51] = 16'sd10;
        fc1_weights[2][52] = 16'sd2;
        fc1_weights[2][53] = 16'sd-17;
        fc1_weights[2][54] = 16'sd-28;
        fc1_weights[2][55] = 16'sd6;
        fc1_weights[2][56] = 16'sd16;
        fc1_weights[2][57] = 16'sd83;
        fc1_weights[2][58] = 16'sd54;
        fc1_weights[2][59] = 16'sd29;
        fc1_weights[2][60] = 16'sd19;
        fc1_weights[2][61] = 16'sd-25;
        fc1_weights[2][62] = 16'sd-79;
        fc1_weights[2][63] = 16'sd-20;
        fc1_weights[2][64] = 16'sd2;
        fc1_weights[2][65] = 16'sd34;
        fc1_weights[2][66] = 16'sd28;
        fc1_weights[2][67] = 16'sd52;
        fc1_weights[2][68] = 16'sd31;
        fc1_weights[2][69] = 16'sd33;
        fc1_weights[2][70] = 16'sd64;
        fc1_weights[2][71] = 16'sd-4;
        fc1_weights[2][72] = 16'sd24;
        fc1_weights[2][73] = 16'sd14;
        fc1_weights[2][74] = 16'sd-39;
        fc1_weights[2][75] = 16'sd-64;
        fc1_weights[2][76] = 16'sd5;
        fc1_weights[2][77] = 16'sd72;
        fc1_weights[2][78] = 16'sd29;
        fc1_weights[2][79] = 16'sd47;
        fc1_weights[2][80] = 16'sd-18;
        fc1_weights[2][81] = 16'sd-52;
        fc1_weights[2][82] = 16'sd-15;
        fc1_weights[2][83] = 16'sd4;
        fc1_weights[2][84] = 16'sd26;
        fc1_weights[2][85] = 16'sd-23;
        fc1_weights[2][86] = 16'sd-31;
        fc1_weights[2][87] = 16'sd-40;
        fc1_weights[2][88] = 16'sd-64;
        fc1_weights[2][89] = 16'sd9;
        fc1_weights[2][90] = 16'sd26;
        fc1_weights[2][91] = 16'sd32;
        fc1_weights[2][92] = 16'sd41;
        fc1_weights[2][93] = 16'sd75;
        fc1_weights[2][94] = 16'sd-21;
        fc1_weights[2][95] = 16'sd46;
        fc1_weights[2][96] = 16'sd45;
        fc1_weights[2][97] = 16'sd81;
        fc1_weights[2][98] = 16'sd43;
        fc1_weights[2][99] = 16'sd-2;
        fc1_weights[2][100] = 16'sd-40;
        fc1_weights[2][101] = 16'sd-45;
        fc1_weights[2][102] = 16'sd-32;
        fc1_weights[2][103] = 16'sd-12;
        fc1_weights[2][104] = 16'sd49;
        fc1_weights[2][105] = 16'sd-34;
        fc1_weights[2][106] = 16'sd26;
        fc1_weights[2][107] = 16'sd-54;
        fc1_weights[2][108] = 16'sd-2;
        fc1_weights[2][109] = 16'sd2;
        fc1_weights[2][110] = 16'sd80;
        fc1_weights[2][111] = 16'sd-32;
        fc1_weights[2][112] = 16'sd7;
        fc1_weights[2][113] = 16'sd-2;
        fc1_weights[2][114] = 16'sd-8;
        fc1_weights[2][115] = 16'sd0;
        fc1_weights[2][116] = 16'sd-45;
        fc1_weights[2][117] = 16'sd13;
        fc1_weights[2][118] = 16'sd-3;
        fc1_weights[2][119] = 16'sd-21;
        fc1_weights[2][120] = 16'sd12;
        fc1_weights[2][121] = 16'sd-75;
        fc1_weights[2][122] = 16'sd-19;
        fc1_weights[2][123] = 16'sd-25;
        fc1_weights[2][124] = 16'sd-103;
        fc1_weights[2][125] = 16'sd-78;
        fc1_weights[2][126] = 16'sd-75;
        fc1_weights[2][127] = 16'sd-4;
        fc1_weights[2][128] = 16'sd-35;
        fc1_weights[2][129] = 16'sd-15;
        fc1_weights[2][130] = 16'sd-33;
        fc1_weights[2][131] = 16'sd-10;
        fc1_weights[2][132] = 16'sd-8;
        fc1_weights[2][133] = 16'sd41;
        fc1_weights[2][134] = 16'sd29;
        fc1_weights[2][135] = 16'sd84;
        fc1_weights[2][136] = 16'sd17;
        fc1_weights[2][137] = 16'sd76;
        fc1_weights[2][138] = 16'sd145;
        fc1_weights[2][139] = 16'sd13;
        fc1_weights[2][140] = 16'sd-13;
        fc1_weights[2][141] = 16'sd-61;
        fc1_weights[2][142] = 16'sd-65;
        fc1_weights[2][143] = 16'sd-43;
        fc1_weights[2][144] = 16'sd76;
        fc1_weights[2][145] = 16'sd-12;
        fc1_weights[2][146] = 16'sd0;
        fc1_weights[2][147] = 16'sd7;
        fc1_weights[2][148] = 16'sd-30;
        fc1_weights[2][149] = 16'sd-13;
        fc1_weights[2][150] = 16'sd-4;
        fc1_weights[2][151] = 16'sd18;
        fc1_weights[2][152] = 16'sd6;
        fc1_weights[2][153] = 16'sd18;
        fc1_weights[2][154] = 16'sd38;
        fc1_weights[2][155] = 16'sd59;
        fc1_weights[2][156] = 16'sd8;
        fc1_weights[2][157] = 16'sd13;
        fc1_weights[2][158] = 16'sd-3;
        fc1_weights[2][159] = 16'sd23;
        fc1_weights[2][160] = 16'sd43;
        fc1_weights[2][161] = 16'sd-14;
        fc1_weights[2][162] = 16'sd-41;
        fc1_weights[2][163] = 16'sd-7;
        fc1_weights[2][164] = 16'sd-57;
        fc1_weights[2][165] = 16'sd26;
        fc1_weights[2][166] = 16'sd19;
        fc1_weights[2][167] = 16'sd-4;
        fc1_weights[2][168] = 16'sd32;
        fc1_weights[2][169] = 16'sd24;
        fc1_weights[2][170] = 16'sd57;
        fc1_weights[2][171] = 16'sd58;
        fc1_weights[2][172] = 16'sd47;
        fc1_weights[2][173] = 16'sd49;
        fc1_weights[2][174] = 16'sd36;
        fc1_weights[2][175] = 16'sd61;
        fc1_weights[2][176] = 16'sd24;
        fc1_weights[2][177] = 16'sd16;
        fc1_weights[2][178] = 16'sd-1;
        fc1_weights[2][179] = 16'sd61;
        fc1_weights[2][180] = 16'sd15;
        fc1_weights[2][181] = 16'sd7;
        fc1_weights[2][182] = 16'sd41;
        fc1_weights[2][183] = 16'sd24;
        fc1_weights[2][184] = 16'sd-19;
        fc1_weights[2][185] = 16'sd-2;
        fc1_weights[2][186] = 16'sd2;
        fc1_weights[2][187] = 16'sd-29;
        fc1_weights[2][188] = 16'sd-24;
        fc1_weights[2][189] = 16'sd-52;
        fc1_weights[2][190] = 16'sd32;
        fc1_weights[2][191] = 16'sd15;
        fc1_weights[2][192] = 16'sd-15;
        fc1_weights[2][193] = 16'sd8;
        fc1_weights[2][194] = 16'sd7;
        fc1_weights[2][195] = 16'sd24;
        fc1_weights[2][196] = 16'sd-13;
        fc1_weights[2][197] = 16'sd47;
        fc1_weights[2][198] = 16'sd66;
        fc1_weights[2][199] = 16'sd48;
        fc1_weights[2][200] = 16'sd20;
        fc1_weights[2][201] = 16'sd-13;
        fc1_weights[2][202] = 16'sd-4;
        fc1_weights[2][203] = 16'sd89;
        fc1_weights[2][204] = 16'sd29;
        fc1_weights[2][205] = 16'sd80;
        fc1_weights[2][206] = 16'sd-19;
        fc1_weights[2][207] = 16'sd-12;
        fc1_weights[3][0] = 16'sd36;
        fc1_weights[3][1] = 16'sd30;
        fc1_weights[3][2] = 16'sd-13;
        fc1_weights[3][3] = 16'sd27;
        fc1_weights[3][4] = 16'sd-37;
        fc1_weights[3][5] = 16'sd-3;
        fc1_weights[3][6] = 16'sd-27;
        fc1_weights[3][7] = 16'sd2;
        fc1_weights[3][8] = 16'sd17;
        fc1_weights[3][9] = 16'sd15;
        fc1_weights[3][10] = 16'sd14;
        fc1_weights[3][11] = 16'sd46;
        fc1_weights[3][12] = 16'sd-25;
        fc1_weights[3][13] = 16'sd14;
        fc1_weights[3][14] = 16'sd-61;
        fc1_weights[3][15] = 16'sd-20;
        fc1_weights[3][16] = 16'sd3;
        fc1_weights[3][17] = 16'sd-11;
        fc1_weights[3][18] = 16'sd15;
        fc1_weights[3][19] = 16'sd74;
        fc1_weights[3][20] = 16'sd91;
        fc1_weights[3][21] = 16'sd54;
        fc1_weights[3][22] = 16'sd5;
        fc1_weights[3][23] = 16'sd24;
        fc1_weights[3][24] = 16'sd44;
        fc1_weights[3][25] = 16'sd-6;
        fc1_weights[3][26] = 16'sd22;
        fc1_weights[3][27] = 16'sd-32;
        fc1_weights[3][28] = 16'sd82;
        fc1_weights[3][29] = 16'sd27;
        fc1_weights[3][30] = 16'sd-5;
        fc1_weights[3][31] = 16'sd-58;
        fc1_weights[3][32] = 16'sd57;
        fc1_weights[3][33] = 16'sd137;
        fc1_weights[3][34] = 16'sd-4;
        fc1_weights[3][35] = 16'sd6;
        fc1_weights[3][36] = 16'sd26;
        fc1_weights[3][37] = 16'sd-58;
        fc1_weights[3][38] = 16'sd-69;
        fc1_weights[3][39] = 16'sd-29;
        fc1_weights[3][40] = 16'sd-3;
        fc1_weights[3][41] = 16'sd-48;
        fc1_weights[3][42] = 16'sd-31;
        fc1_weights[3][43] = 16'sd55;
        fc1_weights[3][44] = 16'sd-3;
        fc1_weights[3][45] = 16'sd79;
        fc1_weights[3][46] = 16'sd102;
        fc1_weights[3][47] = 16'sd88;
        fc1_weights[3][48] = 16'sd2;
        fc1_weights[3][49] = 16'sd-11;
        fc1_weights[3][50] = 16'sd33;
        fc1_weights[3][51] = 16'sd69;
        fc1_weights[3][52] = 16'sd-62;
        fc1_weights[3][53] = 16'sd23;
        fc1_weights[3][54] = 16'sd44;
        fc1_weights[3][55] = 16'sd98;
        fc1_weights[3][56] = 16'sd-22;
        fc1_weights[3][57] = 16'sd-40;
        fc1_weights[3][58] = 16'sd18;
        fc1_weights[3][59] = 16'sd13;
        fc1_weights[3][60] = 16'sd24;
        fc1_weights[3][61] = 16'sd-43;
        fc1_weights[3][62] = 16'sd-6;
        fc1_weights[3][63] = 16'sd-43;
        fc1_weights[3][64] = 16'sd-40;
        fc1_weights[3][65] = 16'sd-10;
        fc1_weights[3][66] = 16'sd12;
        fc1_weights[3][67] = 16'sd-50;
        fc1_weights[3][68] = 16'sd50;
        fc1_weights[3][69] = 16'sd69;
        fc1_weights[3][70] = 16'sd-10;
        fc1_weights[3][71] = 16'sd-2;
        fc1_weights[3][72] = 16'sd47;
        fc1_weights[3][73] = 16'sd-9;
        fc1_weights[3][74] = 16'sd-44;
        fc1_weights[3][75] = 16'sd-12;
        fc1_weights[3][76] = 16'sd-46;
        fc1_weights[3][77] = 16'sd24;
        fc1_weights[3][78] = 16'sd-73;
        fc1_weights[3][79] = 16'sd26;
        fc1_weights[3][80] = 16'sd7;
        fc1_weights[3][81] = 16'sd-22;
        fc1_weights[3][82] = 16'sd18;
        fc1_weights[3][83] = 16'sd-3;
        fc1_weights[3][84] = 16'sd14;
        fc1_weights[3][85] = 16'sd95;
        fc1_weights[3][86] = 16'sd103;
        fc1_weights[3][87] = 16'sd4;
        fc1_weights[3][88] = 16'sd11;
        fc1_weights[3][89] = 16'sd59;
        fc1_weights[3][90] = 16'sd9;
        fc1_weights[3][91] = 16'sd1;
        fc1_weights[3][92] = 16'sd49;
        fc1_weights[3][93] = 16'sd14;
        fc1_weights[3][94] = 16'sd100;
        fc1_weights[3][95] = 16'sd27;
        fc1_weights[3][96] = 16'sd-38;
        fc1_weights[3][97] = 16'sd-79;
        fc1_weights[3][98] = 16'sd-11;
        fc1_weights[3][99] = 16'sd39;
        fc1_weights[3][100] = 16'sd-58;
        fc1_weights[3][101] = 16'sd-15;
        fc1_weights[3][102] = 16'sd112;
        fc1_weights[3][103] = 16'sd41;
        fc1_weights[3][104] = 16'sd-18;
        fc1_weights[3][105] = 16'sd-1;
        fc1_weights[3][106] = 16'sd-8;
        fc1_weights[3][107] = 16'sd24;
        fc1_weights[3][108] = 16'sd-31;
        fc1_weights[3][109] = 16'sd-32;
        fc1_weights[3][110] = 16'sd-15;
        fc1_weights[3][111] = 16'sd-64;
        fc1_weights[3][112] = 16'sd-50;
        fc1_weights[3][113] = 16'sd93;
        fc1_weights[3][114] = 16'sd31;
        fc1_weights[3][115] = 16'sd-30;
        fc1_weights[3][116] = 16'sd13;
        fc1_weights[3][117] = 16'sd57;
        fc1_weights[3][118] = 16'sd-34;
        fc1_weights[3][119] = 16'sd22;
        fc1_weights[3][120] = 16'sd6;
        fc1_weights[3][121] = 16'sd40;
        fc1_weights[3][122] = 16'sd19;
        fc1_weights[3][123] = 16'sd-21;
        fc1_weights[3][124] = 16'sd-30;
        fc1_weights[3][125] = 16'sd30;
        fc1_weights[3][126] = 16'sd-29;
        fc1_weights[3][127] = 16'sd-12;
        fc1_weights[3][128] = 16'sd-91;
        fc1_weights[3][129] = 16'sd-17;
        fc1_weights[3][130] = 16'sd-30;
        fc1_weights[3][131] = 16'sd-85;
        fc1_weights[3][132] = 16'sd-16;
        fc1_weights[3][133] = 16'sd-70;
        fc1_weights[3][134] = 16'sd-2;
        fc1_weights[3][135] = 16'sd10;
        fc1_weights[3][136] = 16'sd-65;
        fc1_weights[3][137] = 16'sd-94;
        fc1_weights[3][138] = 16'sd-105;
        fc1_weights[3][139] = 16'sd47;
        fc1_weights[3][140] = 16'sd-19;
        fc1_weights[3][141] = 16'sd-67;
        fc1_weights[3][142] = 16'sd-86;
        fc1_weights[3][143] = 16'sd-13;
        fc1_weights[3][144] = 16'sd-26;
        fc1_weights[3][145] = 16'sd-50;
        fc1_weights[3][146] = 16'sd-28;
        fc1_weights[3][147] = 16'sd-4;
        fc1_weights[3][148] = 16'sd11;
        fc1_weights[3][149] = 16'sd-20;
        fc1_weights[3][150] = 16'sd-58;
        fc1_weights[3][151] = 16'sd31;
        fc1_weights[3][152] = 16'sd-30;
        fc1_weights[3][153] = 16'sd26;
        fc1_weights[3][154] = 16'sd-3;
        fc1_weights[3][155] = 16'sd51;
        fc1_weights[3][156] = 16'sd25;
        fc1_weights[3][157] = 16'sd36;
        fc1_weights[3][158] = 16'sd19;
        fc1_weights[3][159] = 16'sd44;
        fc1_weights[3][160] = 16'sd-61;
        fc1_weights[3][161] = 16'sd-27;
        fc1_weights[3][162] = 16'sd-65;
        fc1_weights[3][163] = 16'sd-10;
        fc1_weights[3][164] = 16'sd55;
        fc1_weights[3][165] = 16'sd25;
        fc1_weights[3][166] = 16'sd-17;
        fc1_weights[3][167] = 16'sd-8;
        fc1_weights[3][168] = 16'sd-122;
        fc1_weights[3][169] = 16'sd-41;
        fc1_weights[3][170] = 16'sd-52;
        fc1_weights[3][171] = 16'sd10;
        fc1_weights[3][172] = 16'sd-3;
        fc1_weights[3][173] = 16'sd-43;
        fc1_weights[3][174] = 16'sd-19;
        fc1_weights[3][175] = 16'sd9;
        fc1_weights[3][176] = 16'sd37;
        fc1_weights[3][177] = 16'sd44;
        fc1_weights[3][178] = 16'sd9;
        fc1_weights[3][179] = 16'sd2;
        fc1_weights[3][180] = 16'sd3;
        fc1_weights[3][181] = 16'sd8;
        fc1_weights[3][182] = 16'sd-12;
        fc1_weights[3][183] = 16'sd-13;
        fc1_weights[3][184] = 16'sd36;
        fc1_weights[3][185] = 16'sd-3;
        fc1_weights[3][186] = 16'sd-88;
        fc1_weights[3][187] = 16'sd-25;
        fc1_weights[3][188] = 16'sd18;
        fc1_weights[3][189] = 16'sd27;
        fc1_weights[3][190] = 16'sd71;
        fc1_weights[3][191] = 16'sd-16;
        fc1_weights[3][192] = 16'sd-32;
        fc1_weights[3][193] = 16'sd9;
        fc1_weights[3][194] = 16'sd-23;
        fc1_weights[3][195] = 16'sd-5;
        fc1_weights[3][196] = 16'sd-5;
        fc1_weights[3][197] = 16'sd-22;
        fc1_weights[3][198] = 16'sd31;
        fc1_weights[3][199] = 16'sd50;
        fc1_weights[3][200] = 16'sd25;
        fc1_weights[3][201] = 16'sd13;
        fc1_weights[3][202] = 16'sd-48;
        fc1_weights[3][203] = 16'sd2;
        fc1_weights[3][204] = 16'sd3;
        fc1_weights[3][205] = 16'sd-8;
        fc1_weights[3][206] = 16'sd24;
        fc1_weights[3][207] = 16'sd-6;
        fc1_weights[4][0] = 16'sd43;
        fc1_weights[4][1] = 16'sd27;
        fc1_weights[4][2] = 16'sd51;
        fc1_weights[4][3] = 16'sd-22;
        fc1_weights[4][4] = 16'sd23;
        fc1_weights[4][5] = 16'sd12;
        fc1_weights[4][6] = 16'sd8;
        fc1_weights[4][7] = 16'sd-24;
        fc1_weights[4][8] = 16'sd24;
        fc1_weights[4][9] = 16'sd30;
        fc1_weights[4][10] = 16'sd-10;
        fc1_weights[4][11] = 16'sd45;
        fc1_weights[4][12] = 16'sd32;
        fc1_weights[4][13] = 16'sd43;
        fc1_weights[4][14] = 16'sd42;
        fc1_weights[4][15] = 16'sd-50;
        fc1_weights[4][16] = 16'sd-6;
        fc1_weights[4][17] = 16'sd32;
        fc1_weights[4][18] = 16'sd-36;
        fc1_weights[4][19] = 16'sd-37;
        fc1_weights[4][20] = 16'sd-35;
        fc1_weights[4][21] = 16'sd-47;
        fc1_weights[4][22] = 16'sd-17;
        fc1_weights[4][23] = 16'sd17;
        fc1_weights[4][24] = 16'sd-45;
        fc1_weights[4][25] = 16'sd4;
        fc1_weights[4][26] = 16'sd69;
        fc1_weights[4][27] = 16'sd37;
        fc1_weights[4][28] = 16'sd41;
        fc1_weights[4][29] = 16'sd-10;
        fc1_weights[4][30] = 16'sd-12;
        fc1_weights[4][31] = 16'sd5;
        fc1_weights[4][32] = 16'sd40;
        fc1_weights[4][33] = 16'sd-4;
        fc1_weights[4][34] = 16'sd-10;
        fc1_weights[4][35] = 16'sd21;
        fc1_weights[4][36] = 16'sd11;
        fc1_weights[4][37] = 16'sd-3;
        fc1_weights[4][38] = 16'sd76;
        fc1_weights[4][39] = 16'sd50;
        fc1_weights[4][40] = 16'sd-54;
        fc1_weights[4][41] = 16'sd-5;
        fc1_weights[4][42] = 16'sd25;
        fc1_weights[4][43] = 16'sd-51;
        fc1_weights[4][44] = 16'sd-11;
        fc1_weights[4][45] = 16'sd7;
        fc1_weights[4][46] = 16'sd-30;
        fc1_weights[4][47] = 16'sd-25;
        fc1_weights[4][48] = 16'sd-58;
        fc1_weights[4][49] = 16'sd-14;
        fc1_weights[4][50] = 16'sd4;
        fc1_weights[4][51] = 16'sd36;
        fc1_weights[4][52] = 16'sd32;
        fc1_weights[4][53] = 16'sd-16;
        fc1_weights[4][54] = 16'sd-30;
        fc1_weights[4][55] = 16'sd-34;
        fc1_weights[4][56] = 16'sd-53;
        fc1_weights[4][57] = 16'sd-12;
        fc1_weights[4][58] = 16'sd10;
        fc1_weights[4][59] = 16'sd-1;
        fc1_weights[4][60] = 16'sd-16;
        fc1_weights[4][61] = 16'sd-5;
        fc1_weights[4][62] = 16'sd-29;
        fc1_weights[4][63] = 16'sd63;
        fc1_weights[4][64] = 16'sd-24;
        fc1_weights[4][65] = 16'sd-38;
        fc1_weights[4][66] = 16'sd-21;
        fc1_weights[4][67] = 16'sd-51;
        fc1_weights[4][68] = 16'sd29;
        fc1_weights[4][69] = 16'sd40;
        fc1_weights[4][70] = 16'sd58;
        fc1_weights[4][71] = 16'sd66;
        fc1_weights[4][72] = 16'sd-41;
        fc1_weights[4][73] = 16'sd29;
        fc1_weights[4][74] = 16'sd4;
        fc1_weights[4][75] = 16'sd2;
        fc1_weights[4][76] = 16'sd-40;
        fc1_weights[4][77] = 16'sd-5;
        fc1_weights[4][78] = 16'sd-11;
        fc1_weights[4][79] = 16'sd-36;
        fc1_weights[4][80] = 16'sd-18;
        fc1_weights[4][81] = 16'sd-52;
        fc1_weights[4][82] = 16'sd-64;
        fc1_weights[4][83] = 16'sd-7;
        fc1_weights[4][84] = 16'sd-29;
        fc1_weights[4][85] = 16'sd-18;
        fc1_weights[4][86] = 16'sd-41;
        fc1_weights[4][87] = 16'sd-53;
        fc1_weights[4][88] = 16'sd5;
        fc1_weights[4][89] = 16'sd-82;
        fc1_weights[4][90] = 16'sd5;
        fc1_weights[4][91] = 16'sd-80;
        fc1_weights[4][92] = 16'sd-22;
        fc1_weights[4][93] = 16'sd-49;
        fc1_weights[4][94] = 16'sd-28;
        fc1_weights[4][95] = 16'sd49;
        fc1_weights[4][96] = 16'sd43;
        fc1_weights[4][97] = 16'sd46;
        fc1_weights[4][98] = 16'sd-16;
        fc1_weights[4][99] = 16'sd-38;
        fc1_weights[4][100] = 16'sd-30;
        fc1_weights[4][101] = 16'sd-66;
        fc1_weights[4][102] = 16'sd-40;
        fc1_weights[4][103] = 16'sd11;
        fc1_weights[4][104] = 16'sd-29;
        fc1_weights[4][105] = 16'sd0;
        fc1_weights[4][106] = 16'sd-4;
        fc1_weights[4][107] = 16'sd-7;
        fc1_weights[4][108] = 16'sd-35;
        fc1_weights[4][109] = 16'sd-7;
        fc1_weights[4][110] = 16'sd-39;
        fc1_weights[4][111] = 16'sd-38;
        fc1_weights[4][112] = 16'sd18;
        fc1_weights[4][113] = 16'sd-4;
        fc1_weights[4][114] = 16'sd-59;
        fc1_weights[4][115] = 16'sd-55;
        fc1_weights[4][116] = 16'sd-21;
        fc1_weights[4][117] = 16'sd-67;
        fc1_weights[4][118] = 16'sd-33;
        fc1_weights[4][119] = 16'sd-33;
        fc1_weights[4][120] = 16'sd45;
        fc1_weights[4][121] = 16'sd14;
        fc1_weights[4][122] = 16'sd22;
        fc1_weights[4][123] = 16'sd26;
        fc1_weights[4][124] = 16'sd44;
        fc1_weights[4][125] = 16'sd-18;
        fc1_weights[4][126] = 16'sd-19;
        fc1_weights[4][127] = 16'sd1;
        fc1_weights[4][128] = 16'sd10;
        fc1_weights[4][129] = 16'sd43;
        fc1_weights[4][130] = 16'sd-24;
        fc1_weights[4][131] = 16'sd-8;
        fc1_weights[4][132] = 16'sd-22;
        fc1_weights[4][133] = 16'sd-12;
        fc1_weights[4][134] = 16'sd-37;
        fc1_weights[4][135] = 16'sd-50;
        fc1_weights[4][136] = 16'sd-37;
        fc1_weights[4][137] = 16'sd-31;
        fc1_weights[4][138] = 16'sd9;
        fc1_weights[4][139] = 16'sd17;
        fc1_weights[4][140] = 16'sd-15;
        fc1_weights[4][141] = 16'sd-5;
        fc1_weights[4][142] = 16'sd6;
        fc1_weights[4][143] = 16'sd-64;
        fc1_weights[4][144] = 16'sd1;
        fc1_weights[4][145] = 16'sd-23;
        fc1_weights[4][146] = 16'sd-34;
        fc1_weights[4][147] = 16'sd6;
        fc1_weights[4][148] = 16'sd8;
        fc1_weights[4][149] = 16'sd8;
        fc1_weights[4][150] = 16'sd20;
        fc1_weights[4][151] = 16'sd-19;
        fc1_weights[4][152] = 16'sd-33;
        fc1_weights[4][153] = 16'sd-34;
        fc1_weights[4][154] = 16'sd12;
        fc1_weights[4][155] = 16'sd20;
        fc1_weights[4][156] = 16'sd-26;
        fc1_weights[4][157] = 16'sd-13;
        fc1_weights[4][158] = 16'sd-22;
        fc1_weights[4][159] = 16'sd-24;
        fc1_weights[4][160] = 16'sd33;
        fc1_weights[4][161] = 16'sd47;
        fc1_weights[4][162] = 16'sd-2;
        fc1_weights[4][163] = 16'sd35;
        fc1_weights[4][164] = 16'sd12;
        fc1_weights[4][165] = 16'sd31;
        fc1_weights[4][166] = 16'sd-48;
        fc1_weights[4][167] = 16'sd-21;
        fc1_weights[4][168] = 16'sd-61;
        fc1_weights[4][169] = 16'sd-20;
        fc1_weights[4][170] = 16'sd25;
        fc1_weights[4][171] = 16'sd-9;
        fc1_weights[4][172] = 16'sd-17;
        fc1_weights[4][173] = 16'sd-10;
        fc1_weights[4][174] = 16'sd-5;
        fc1_weights[4][175] = 16'sd-18;
        fc1_weights[4][176] = 16'sd-13;
        fc1_weights[4][177] = 16'sd27;
        fc1_weights[4][178] = 16'sd-13;
        fc1_weights[4][179] = 16'sd-50;
        fc1_weights[4][180] = 16'sd-5;
        fc1_weights[4][181] = 16'sd-31;
        fc1_weights[4][182] = 16'sd-10;
        fc1_weights[4][183] = 16'sd-38;
        fc1_weights[4][184] = 16'sd12;
        fc1_weights[4][185] = 16'sd-32;
        fc1_weights[4][186] = 16'sd10;
        fc1_weights[4][187] = 16'sd19;
        fc1_weights[4][188] = 16'sd-24;
        fc1_weights[4][189] = 16'sd27;
        fc1_weights[4][190] = 16'sd37;
        fc1_weights[4][191] = 16'sd-47;
        fc1_weights[4][192] = 16'sd3;
        fc1_weights[4][193] = 16'sd-37;
        fc1_weights[4][194] = 16'sd20;
        fc1_weights[4][195] = 16'sd5;
        fc1_weights[4][196] = 16'sd42;
        fc1_weights[4][197] = 16'sd-34;
        fc1_weights[4][198] = 16'sd9;
        fc1_weights[4][199] = 16'sd21;
        fc1_weights[4][200] = 16'sd5;
        fc1_weights[4][201] = 16'sd17;
        fc1_weights[4][202] = 16'sd-22;
        fc1_weights[4][203] = 16'sd28;
        fc1_weights[4][204] = 16'sd-22;
        fc1_weights[4][205] = 16'sd9;
        fc1_weights[4][206] = 16'sd30;
        fc1_weights[4][207] = 16'sd6;
        fc1_weights[5][0] = 16'sd-45;
        fc1_weights[5][1] = 16'sd-16;
        fc1_weights[5][2] = 16'sd20;
        fc1_weights[5][3] = 16'sd40;
        fc1_weights[5][4] = 16'sd51;
        fc1_weights[5][5] = 16'sd17;
        fc1_weights[5][6] = 16'sd5;
        fc1_weights[5][7] = 16'sd45;
        fc1_weights[5][8] = 16'sd10;
        fc1_weights[5][9] = 16'sd4;
        fc1_weights[5][10] = 16'sd-23;
        fc1_weights[5][11] = 16'sd22;
        fc1_weights[5][12] = 16'sd50;
        fc1_weights[5][13] = 16'sd50;
        fc1_weights[5][14] = 16'sd50;
        fc1_weights[5][15] = 16'sd-15;
        fc1_weights[5][16] = 16'sd1;
        fc1_weights[5][17] = 16'sd53;
        fc1_weights[5][18] = 16'sd35;
        fc1_weights[5][19] = 16'sd22;
        fc1_weights[5][20] = 16'sd45;
        fc1_weights[5][21] = 16'sd49;
        fc1_weights[5][22] = 16'sd58;
        fc1_weights[5][23] = 16'sd64;
        fc1_weights[5][24] = 16'sd48;
        fc1_weights[5][25] = 16'sd25;
        fc1_weights[5][26] = 16'sd-3;
        fc1_weights[5][27] = 16'sd-10;
        fc1_weights[5][28] = 16'sd6;
        fc1_weights[5][29] = 16'sd45;
        fc1_weights[5][30] = 16'sd-1;
        fc1_weights[5][31] = 16'sd-4;
        fc1_weights[5][32] = 16'sd3;
        fc1_weights[5][33] = 16'sd15;
        fc1_weights[5][34] = 16'sd30;
        fc1_weights[5][35] = 16'sd1;
        fc1_weights[5][36] = 16'sd-25;
        fc1_weights[5][37] = 16'sd-11;
        fc1_weights[5][38] = 16'sd24;
        fc1_weights[5][39] = 16'sd65;
        fc1_weights[5][40] = 16'sd-20;
        fc1_weights[5][41] = 16'sd16;
        fc1_weights[5][42] = 16'sd37;
        fc1_weights[5][43] = 16'sd-47;
        fc1_weights[5][44] = 16'sd18;
        fc1_weights[5][45] = 16'sd14;
        fc1_weights[5][46] = 16'sd43;
        fc1_weights[5][47] = 16'sd28;
        fc1_weights[5][48] = 16'sd37;
        fc1_weights[5][49] = 16'sd-3;
        fc1_weights[5][50] = 16'sd29;
        fc1_weights[5][51] = 16'sd9;
        fc1_weights[5][52] = 16'sd-27;
        fc1_weights[5][53] = 16'sd-43;
        fc1_weights[5][54] = 16'sd-73;
        fc1_weights[5][55] = 16'sd-41;
        fc1_weights[5][56] = 16'sd-42;
        fc1_weights[5][57] = 16'sd-31;
        fc1_weights[5][58] = 16'sd-3;
        fc1_weights[5][59] = 16'sd20;
        fc1_weights[5][60] = 16'sd-6;
        fc1_weights[5][61] = 16'sd12;
        fc1_weights[5][62] = 16'sd16;
        fc1_weights[5][63] = 16'sd-2;
        fc1_weights[5][64] = 16'sd0;
        fc1_weights[5][65] = 16'sd0;
        fc1_weights[5][66] = 16'sd18;
        fc1_weights[5][67] = 16'sd-31;
        fc1_weights[5][68] = 16'sd-5;
        fc1_weights[5][69] = 16'sd-28;
        fc1_weights[5][70] = 16'sd3;
        fc1_weights[5][71] = 16'sd5;
        fc1_weights[5][72] = 16'sd26;
        fc1_weights[5][73] = 16'sd48;
        fc1_weights[5][74] = 16'sd40;
        fc1_weights[5][75] = 16'sd14;
        fc1_weights[5][76] = 16'sd-27;
        fc1_weights[5][77] = 16'sd-21;
        fc1_weights[5][78] = 16'sd-44;
        fc1_weights[5][79] = 16'sd-27;
        fc1_weights[5][80] = 16'sd-26;
        fc1_weights[5][81] = 16'sd-20;
        fc1_weights[5][82] = 16'sd-43;
        fc1_weights[5][83] = 16'sd14;
        fc1_weights[5][84] = 16'sd14;
        fc1_weights[5][85] = 16'sd16;
        fc1_weights[5][86] = 16'sd25;
        fc1_weights[5][87] = 16'sd24;
        fc1_weights[5][88] = 16'sd31;
        fc1_weights[5][89] = 16'sd-14;
        fc1_weights[5][90] = 16'sd19;
        fc1_weights[5][91] = 16'sd-25;
        fc1_weights[5][92] = 16'sd24;
        fc1_weights[5][93] = 16'sd-89;
        fc1_weights[5][94] = 16'sd-52;
        fc1_weights[5][95] = 16'sd-33;
        fc1_weights[5][96] = 16'sd21;
        fc1_weights[5][97] = 16'sd-61;
        fc1_weights[5][98] = 16'sd3;
        fc1_weights[5][99] = 16'sd-22;
        fc1_weights[5][100] = 16'sd7;
        fc1_weights[5][101] = 16'sd5;
        fc1_weights[5][102] = 16'sd-11;
        fc1_weights[5][103] = 16'sd-9;
        fc1_weights[5][104] = 16'sd0;
        fc1_weights[5][105] = 16'sd-18;
        fc1_weights[5][106] = 16'sd9;
        fc1_weights[5][107] = 16'sd-3;
        fc1_weights[5][108] = 16'sd3;
        fc1_weights[5][109] = 16'sd36;
        fc1_weights[5][110] = 16'sd67;
        fc1_weights[5][111] = 16'sd72;
        fc1_weights[5][112] = 16'sd-17;
        fc1_weights[5][113] = 16'sd-75;
        fc1_weights[5][114] = 16'sd18;
        fc1_weights[5][115] = 16'sd36;
        fc1_weights[5][116] = 16'sd17;
        fc1_weights[5][117] = 16'sd-14;
        fc1_weights[5][118] = 16'sd18;
        fc1_weights[5][119] = 16'sd-17;
        fc1_weights[5][120] = 16'sd-38;
        fc1_weights[5][121] = 16'sd7;
        fc1_weights[5][122] = 16'sd18;
        fc1_weights[5][123] = 16'sd-59;
        fc1_weights[5][124] = 16'sd43;
        fc1_weights[5][125] = 16'sd-8;
        fc1_weights[5][126] = 16'sd42;
        fc1_weights[5][127] = 16'sd-11;
        fc1_weights[5][128] = 16'sd66;
        fc1_weights[5][129] = 16'sd32;
        fc1_weights[5][130] = 16'sd35;
        fc1_weights[5][131] = 16'sd32;
        fc1_weights[5][132] = 16'sd1;
        fc1_weights[5][133] = 16'sd-28;
        fc1_weights[5][134] = 16'sd-11;
        fc1_weights[5][135] = 16'sd-47;
        fc1_weights[5][136] = 16'sd3;
        fc1_weights[5][137] = 16'sd23;
        fc1_weights[5][138] = 16'sd-24;
        fc1_weights[5][139] = 16'sd-41;
        fc1_weights[5][140] = 16'sd9;
        fc1_weights[5][141] = 16'sd90;
        fc1_weights[5][142] = 16'sd16;
        fc1_weights[5][143] = 16'sd1;
        fc1_weights[5][144] = 16'sd18;
        fc1_weights[5][145] = 16'sd83;
        fc1_weights[5][146] = 16'sd9;
        fc1_weights[5][147] = 16'sd24;
        fc1_weights[5][148] = 16'sd-26;
        fc1_weights[5][149] = 16'sd-16;
        fc1_weights[5][150] = 16'sd5;
        fc1_weights[5][151] = 16'sd-23;
        fc1_weights[5][152] = 16'sd23;
        fc1_weights[5][153] = 16'sd4;
        fc1_weights[5][154] = 16'sd28;
        fc1_weights[5][155] = 16'sd-28;
        fc1_weights[5][156] = 16'sd-6;
        fc1_weights[5][157] = 16'sd-12;
        fc1_weights[5][158] = 16'sd1;
        fc1_weights[5][159] = 16'sd-2;
        fc1_weights[5][160] = 16'sd-5;
        fc1_weights[5][161] = 16'sd38;
        fc1_weights[5][162] = 16'sd-28;
        fc1_weights[5][163] = 16'sd-8;
        fc1_weights[5][164] = 16'sd-15;
        fc1_weights[5][165] = 16'sd-62;
        fc1_weights[5][166] = 16'sd-3;
        fc1_weights[5][167] = 16'sd-19;
        fc1_weights[5][168] = 16'sd-10;
        fc1_weights[5][169] = 16'sd3;
        fc1_weights[5][170] = 16'sd24;
        fc1_weights[5][171] = 16'sd27;
        fc1_weights[5][172] = 16'sd21;
        fc1_weights[5][173] = 16'sd5;
        fc1_weights[5][174] = 16'sd9;
        fc1_weights[5][175] = 16'sd-10;
        fc1_weights[5][176] = 16'sd-47;
        fc1_weights[5][177] = 16'sd-17;
        fc1_weights[5][178] = 16'sd45;
        fc1_weights[5][179] = 16'sd-53;
        fc1_weights[5][180] = 16'sd-37;
        fc1_weights[5][181] = 16'sd-13;
        fc1_weights[5][182] = 16'sd-25;
        fc1_weights[5][183] = 16'sd-34;
        fc1_weights[5][184] = 16'sd-16;
        fc1_weights[5][185] = 16'sd-39;
        fc1_weights[5][186] = 16'sd-18;
        fc1_weights[5][187] = 16'sd-26;
        fc1_weights[5][188] = 16'sd-24;
        fc1_weights[5][189] = 16'sd-2;
        fc1_weights[5][190] = 16'sd-76;
        fc1_weights[5][191] = 16'sd-38;
        fc1_weights[5][192] = 16'sd9;
        fc1_weights[5][193] = 16'sd-6;
        fc1_weights[5][194] = 16'sd-24;
        fc1_weights[5][195] = 16'sd3;
        fc1_weights[5][196] = 16'sd-12;
        fc1_weights[5][197] = 16'sd-41;
        fc1_weights[5][198] = 16'sd2;
        fc1_weights[5][199] = 16'sd-2;
        fc1_weights[5][200] = 16'sd45;
        fc1_weights[5][201] = 16'sd18;
        fc1_weights[5][202] = 16'sd75;
        fc1_weights[5][203] = 16'sd-8;
        fc1_weights[5][204] = 16'sd-14;
        fc1_weights[5][205] = 16'sd4;
        fc1_weights[5][206] = 16'sd51;
        fc1_weights[5][207] = 16'sd48;
        fc1_weights[6][0] = 16'sd-5;
        fc1_weights[6][1] = 16'sd-8;
        fc1_weights[6][2] = 16'sd-1;
        fc1_weights[6][3] = 16'sd-23;
        fc1_weights[6][4] = 16'sd41;
        fc1_weights[6][5] = 16'sd5;
        fc1_weights[6][6] = 16'sd-24;
        fc1_weights[6][7] = 16'sd-73;
        fc1_weights[6][8] = 16'sd-9;
        fc1_weights[6][9] = 16'sd6;
        fc1_weights[6][10] = 16'sd-68;
        fc1_weights[6][11] = 16'sd37;
        fc1_weights[6][12] = 16'sd52;
        fc1_weights[6][13] = 16'sd53;
        fc1_weights[6][14] = 16'sd45;
        fc1_weights[6][15] = 16'sd-60;
        fc1_weights[6][16] = 16'sd-14;
        fc1_weights[6][17] = 16'sd54;
        fc1_weights[6][18] = 16'sd-8;
        fc1_weights[6][19] = 16'sd-41;
        fc1_weights[6][20] = 16'sd38;
        fc1_weights[6][21] = 16'sd-30;
        fc1_weights[6][22] = 16'sd-42;
        fc1_weights[6][23] = 16'sd18;
        fc1_weights[6][24] = 16'sd-19;
        fc1_weights[6][25] = 16'sd-37;
        fc1_weights[6][26] = 16'sd7;
        fc1_weights[6][27] = 16'sd20;
        fc1_weights[6][28] = 16'sd-4;
        fc1_weights[6][29] = 16'sd-27;
        fc1_weights[6][30] = 16'sd-10;
        fc1_weights[6][31] = 16'sd20;
        fc1_weights[6][32] = 16'sd-12;
        fc1_weights[6][33] = 16'sd10;
        fc1_weights[6][34] = 16'sd-24;
        fc1_weights[6][35] = 16'sd-30;
        fc1_weights[6][36] = 16'sd-60;
        fc1_weights[6][37] = 16'sd-67;
        fc1_weights[6][38] = 16'sd14;
        fc1_weights[6][39] = 16'sd63;
        fc1_weights[6][40] = 16'sd-133;
        fc1_weights[6][41] = 16'sd-17;
        fc1_weights[6][42] = 16'sd42;
        fc1_weights[6][43] = 16'sd-3;
        fc1_weights[6][44] = 16'sd-17;
        fc1_weights[6][45] = 16'sd11;
        fc1_weights[6][46] = 16'sd24;
        fc1_weights[6][47] = 16'sd54;
        fc1_weights[6][48] = 16'sd-53;
        fc1_weights[6][49] = 16'sd-46;
        fc1_weights[6][50] = 16'sd20;
        fc1_weights[6][51] = 16'sd52;
        fc1_weights[6][52] = 16'sd15;
        fc1_weights[6][53] = 16'sd-37;
        fc1_weights[6][54] = 16'sd-36;
        fc1_weights[6][55] = 16'sd-43;
        fc1_weights[6][56] = 16'sd-54;
        fc1_weights[6][57] = 16'sd-17;
        fc1_weights[6][58] = 16'sd-19;
        fc1_weights[6][59] = 16'sd-13;
        fc1_weights[6][60] = 16'sd-80;
        fc1_weights[6][61] = 16'sd-36;
        fc1_weights[6][62] = 16'sd11;
        fc1_weights[6][63] = 16'sd-41;
        fc1_weights[6][64] = 16'sd-14;
        fc1_weights[6][65] = 16'sd35;
        fc1_weights[6][66] = 16'sd-2;
        fc1_weights[6][67] = 16'sd-19;
        fc1_weights[6][68] = 16'sd-11;
        fc1_weights[6][69] = 16'sd-61;
        fc1_weights[6][70] = 16'sd10;
        fc1_weights[6][71] = 16'sd48;
        fc1_weights[6][72] = 16'sd12;
        fc1_weights[6][73] = 16'sd39;
        fc1_weights[6][74] = 16'sd36;
        fc1_weights[6][75] = 16'sd33;
        fc1_weights[6][76] = 16'sd-31;
        fc1_weights[6][77] = 16'sd10;
        fc1_weights[6][78] = 16'sd-25;
        fc1_weights[6][79] = 16'sd-54;
        fc1_weights[6][80] = 16'sd-21;
        fc1_weights[6][81] = 16'sd-17;
        fc1_weights[6][82] = 16'sd-47;
        fc1_weights[6][83] = 16'sd0;
        fc1_weights[6][84] = 16'sd-10;
        fc1_weights[6][85] = 16'sd28;
        fc1_weights[6][86] = 16'sd-20;
        fc1_weights[6][87] = 16'sd-46;
        fc1_weights[6][88] = 16'sd35;
        fc1_weights[6][89] = 16'sd-84;
        fc1_weights[6][90] = 16'sd-29;
        fc1_weights[6][91] = 16'sd-2;
        fc1_weights[6][92] = 16'sd-11;
        fc1_weights[6][93] = 16'sd-13;
        fc1_weights[6][94] = 16'sd-9;
        fc1_weights[6][95] = 16'sd43;
        fc1_weights[6][96] = 16'sd56;
        fc1_weights[6][97] = 16'sd56;
        fc1_weights[6][98] = 16'sd37;
        fc1_weights[6][99] = 16'sd18;
        fc1_weights[6][100] = 16'sd21;
        fc1_weights[6][101] = 16'sd10;
        fc1_weights[6][102] = 16'sd42;
        fc1_weights[6][103] = 16'sd71;
        fc1_weights[6][104] = 16'sd-25;
        fc1_weights[6][105] = 16'sd-2;
        fc1_weights[6][106] = 16'sd-6;
        fc1_weights[6][107] = 16'sd3;
        fc1_weights[6][108] = 16'sd10;
        fc1_weights[6][109] = 16'sd-13;
        fc1_weights[6][110] = 16'sd-15;
        fc1_weights[6][111] = 16'sd16;
        fc1_weights[6][112] = 16'sd-59;
        fc1_weights[6][113] = 16'sd-38;
        fc1_weights[6][114] = 16'sd-72;
        fc1_weights[6][115] = 16'sd-38;
        fc1_weights[6][116] = 16'sd-23;
        fc1_weights[6][117] = 16'sd-5;
        fc1_weights[6][118] = 16'sd-19;
        fc1_weights[6][119] = 16'sd59;
        fc1_weights[6][120] = 16'sd65;
        fc1_weights[6][121] = 16'sd62;
        fc1_weights[6][122] = 16'sd35;
        fc1_weights[6][123] = 16'sd35;
        fc1_weights[6][124] = 16'sd80;
        fc1_weights[6][125] = 16'sd69;
        fc1_weights[6][126] = 16'sd103;
        fc1_weights[6][127] = 16'sd21;
        fc1_weights[6][128] = 16'sd48;
        fc1_weights[6][129] = 16'sd54;
        fc1_weights[6][130] = 16'sd-26;
        fc1_weights[6][131] = 16'sd-21;
        fc1_weights[6][132] = 16'sd1;
        fc1_weights[6][133] = 16'sd-11;
        fc1_weights[6][134] = 16'sd-6;
        fc1_weights[6][135] = 16'sd-22;
        fc1_weights[6][136] = 16'sd-14;
        fc1_weights[6][137] = 16'sd7;
        fc1_weights[6][138] = 16'sd-39;
        fc1_weights[6][139] = 16'sd14;
        fc1_weights[6][140] = 16'sd10;
        fc1_weights[6][141] = 16'sd34;
        fc1_weights[6][142] = 16'sd12;
        fc1_weights[6][143] = 16'sd24;
        fc1_weights[6][144] = 16'sd-10;
        fc1_weights[6][145] = 16'sd13;
        fc1_weights[6][146] = 16'sd2;
        fc1_weights[6][147] = 16'sd52;
        fc1_weights[6][148] = 16'sd33;
        fc1_weights[6][149] = 16'sd71;
        fc1_weights[6][150] = 16'sd38;
        fc1_weights[6][151] = 16'sd53;
        fc1_weights[6][152] = 16'sd18;
        fc1_weights[6][153] = 16'sd-7;
        fc1_weights[6][154] = 16'sd35;
        fc1_weights[6][155] = 16'sd24;
        fc1_weights[6][156] = 16'sd26;
        fc1_weights[6][157] = 16'sd18;
        fc1_weights[6][158] = 16'sd10;
        fc1_weights[6][159] = 16'sd0;
        fc1_weights[6][160] = 16'sd-11;
        fc1_weights[6][161] = 16'sd50;
        fc1_weights[6][162] = 16'sd-40;
        fc1_weights[6][163] = 16'sd6;
        fc1_weights[6][164] = 16'sd-32;
        fc1_weights[6][165] = 16'sd-37;
        fc1_weights[6][166] = 16'sd-39;
        fc1_weights[6][167] = 16'sd-49;
        fc1_weights[6][168] = 16'sd-38;
        fc1_weights[6][169] = 16'sd14;
        fc1_weights[6][170] = 16'sd50;
        fc1_weights[6][171] = 16'sd10;
        fc1_weights[6][172] = 16'sd-42;
        fc1_weights[6][173] = 16'sd25;
        fc1_weights[6][174] = 16'sd10;
        fc1_weights[6][175] = 16'sd61;
        fc1_weights[6][176] = 16'sd25;
        fc1_weights[6][177] = 16'sd0;
        fc1_weights[6][178] = 16'sd53;
        fc1_weights[6][179] = 16'sd-14;
        fc1_weights[6][180] = 16'sd43;
        fc1_weights[6][181] = 16'sd-11;
        fc1_weights[6][182] = 16'sd-12;
        fc1_weights[6][183] = 16'sd-45;
        fc1_weights[6][184] = 16'sd2;
        fc1_weights[6][185] = 16'sd-23;
        fc1_weights[6][186] = 16'sd-35;
        fc1_weights[6][187] = 16'sd-36;
        fc1_weights[6][188] = 16'sd-58;
        fc1_weights[6][189] = 16'sd3;
        fc1_weights[6][190] = 16'sd12;
        fc1_weights[6][191] = 16'sd-73;
        fc1_weights[6][192] = 16'sd-4;
        fc1_weights[6][193] = 16'sd-42;
        fc1_weights[6][194] = 16'sd9;
        fc1_weights[6][195] = 16'sd7;
        fc1_weights[6][196] = 16'sd62;
        fc1_weights[6][197] = 16'sd-10;
        fc1_weights[6][198] = 16'sd-1;
        fc1_weights[6][199] = 16'sd-4;
        fc1_weights[6][200] = 16'sd-3;
        fc1_weights[6][201] = 16'sd-5;
        fc1_weights[6][202] = 16'sd19;
        fc1_weights[6][203] = 16'sd-20;
        fc1_weights[6][204] = 16'sd-39;
        fc1_weights[6][205] = 16'sd-22;
        fc1_weights[6][206] = 16'sd47;
        fc1_weights[6][207] = 16'sd14;
        fc1_weights[7][0] = 16'sd-8;
        fc1_weights[7][1] = 16'sd4;
        fc1_weights[7][2] = 16'sd-5;
        fc1_weights[7][3] = 16'sd31;
        fc1_weights[7][4] = 16'sd12;
        fc1_weights[7][5] = 16'sd3;
        fc1_weights[7][6] = 16'sd29;
        fc1_weights[7][7] = 16'sd30;
        fc1_weights[7][8] = 16'sd2;
        fc1_weights[7][9] = 16'sd-22;
        fc1_weights[7][10] = 16'sd9;
        fc1_weights[7][11] = 16'sd1;
        fc1_weights[7][12] = 16'sd32;
        fc1_weights[7][13] = 16'sd27;
        fc1_weights[7][14] = 16'sd26;
        fc1_weights[7][15] = 16'sd19;
        fc1_weights[7][16] = 16'sd6;
        fc1_weights[7][17] = 16'sd-6;
        fc1_weights[7][18] = 16'sd-16;
        fc1_weights[7][19] = 16'sd-3;
        fc1_weights[7][20] = 16'sd-12;
        fc1_weights[7][21] = 16'sd-1;
        fc1_weights[7][22] = 16'sd11;
        fc1_weights[7][23] = 16'sd-24;
        fc1_weights[7][24] = 16'sd-7;
        fc1_weights[7][25] = 16'sd0;
        fc1_weights[7][26] = 16'sd10;
        fc1_weights[7][27] = 16'sd-36;
        fc1_weights[7][28] = 16'sd-1;
        fc1_weights[7][29] = 16'sd4;
        fc1_weights[7][30] = 16'sd-7;
        fc1_weights[7][31] = 16'sd-18;
        fc1_weights[7][32] = 16'sd-1;
        fc1_weights[7][33] = 16'sd52;
        fc1_weights[7][34] = 16'sd6;
        fc1_weights[7][35] = 16'sd-1;
        fc1_weights[7][36] = 16'sd25;
        fc1_weights[7][37] = 16'sd33;
        fc1_weights[7][38] = 16'sd-24;
        fc1_weights[7][39] = 16'sd-4;
        fc1_weights[7][40] = 16'sd4;
        fc1_weights[7][41] = 16'sd-15;
        fc1_weights[7][42] = 16'sd-7;
        fc1_weights[7][43] = 16'sd1;
        fc1_weights[7][44] = 16'sd-15;
        fc1_weights[7][45] = 16'sd5;
        fc1_weights[7][46] = 16'sd-7;
        fc1_weights[7][47] = 16'sd-4;
        fc1_weights[7][48] = 16'sd-20;
        fc1_weights[7][49] = 16'sd0;
        fc1_weights[7][50] = 16'sd-14;
        fc1_weights[7][51] = 16'sd-14;
        fc1_weights[7][52] = 16'sd-3;
        fc1_weights[7][53] = 16'sd-18;
        fc1_weights[7][54] = 16'sd-5;
        fc1_weights[7][55] = 16'sd19;
        fc1_weights[7][56] = 16'sd2;
        fc1_weights[7][57] = 16'sd-2;
        fc1_weights[7][58] = 16'sd-29;
        fc1_weights[7][59] = 16'sd-2;
        fc1_weights[7][60] = 16'sd-14;
        fc1_weights[7][61] = 16'sd-12;
        fc1_weights[7][62] = 16'sd15;
        fc1_weights[7][63] = 16'sd4;
        fc1_weights[7][64] = 16'sd-4;
        fc1_weights[7][65] = 16'sd8;
        fc1_weights[7][66] = 16'sd6;
        fc1_weights[7][67] = 16'sd-29;
        fc1_weights[7][68] = 16'sd3;
        fc1_weights[7][69] = 16'sd19;
        fc1_weights[7][70] = 16'sd13;
        fc1_weights[7][71] = 16'sd-14;
        fc1_weights[7][72] = 16'sd8;
        fc1_weights[7][73] = 16'sd-9;
        fc1_weights[7][74] = 16'sd5;
        fc1_weights[7][75] = 16'sd-4;
        fc1_weights[7][76] = 16'sd-27;
        fc1_weights[7][77] = 16'sd4;
        fc1_weights[7][78] = 16'sd11;
        fc1_weights[7][79] = 16'sd29;
        fc1_weights[7][80] = 16'sd11;
        fc1_weights[7][81] = 16'sd0;
        fc1_weights[7][82] = 16'sd6;
        fc1_weights[7][83] = 16'sd-11;
        fc1_weights[7][84] = 16'sd-13;
        fc1_weights[7][85] = 16'sd15;
        fc1_weights[7][86] = 16'sd-17;
        fc1_weights[7][87] = 16'sd5;
        fc1_weights[7][88] = 16'sd13;
        fc1_weights[7][89] = 16'sd15;
        fc1_weights[7][90] = 16'sd-31;
        fc1_weights[7][91] = 16'sd-24;
        fc1_weights[7][92] = 16'sd-29;
        fc1_weights[7][93] = 16'sd3;
        fc1_weights[7][94] = 16'sd-2;
        fc1_weights[7][95] = 16'sd-6;
        fc1_weights[7][96] = 16'sd12;
        fc1_weights[7][97] = 16'sd-1;
        fc1_weights[7][98] = 16'sd-5;
        fc1_weights[7][99] = 16'sd-15;
        fc1_weights[7][100] = 16'sd-17;
        fc1_weights[7][101] = 16'sd-5;
        fc1_weights[7][102] = 16'sd4;
        fc1_weights[7][103] = 16'sd-1;
        fc1_weights[7][104] = 16'sd28;
        fc1_weights[7][105] = 16'sd28;
        fc1_weights[7][106] = 16'sd20;
        fc1_weights[7][107] = 16'sd-17;
        fc1_weights[7][108] = 16'sd-8;
        fc1_weights[7][109] = 16'sd-4;
        fc1_weights[7][110] = 16'sd-21;
        fc1_weights[7][111] = 16'sd-1;
        fc1_weights[7][112] = 16'sd-11;
        fc1_weights[7][113] = 16'sd-18;
        fc1_weights[7][114] = 16'sd44;
        fc1_weights[7][115] = 16'sd28;
        fc1_weights[7][116] = 16'sd4;
        fc1_weights[7][117] = 16'sd-24;
        fc1_weights[7][118] = 16'sd-44;
        fc1_weights[7][119] = 16'sd-41;
        fc1_weights[7][120] = 16'sd-44;
        fc1_weights[7][121] = 16'sd-11;
        fc1_weights[7][122] = 16'sd-10;
        fc1_weights[7][123] = 16'sd-33;
        fc1_weights[7][124] = 16'sd-14;
        fc1_weights[7][125] = 16'sd-15;
        fc1_weights[7][126] = 16'sd-13;
        fc1_weights[7][127] = 16'sd-42;
        fc1_weights[7][128] = 16'sd-37;
        fc1_weights[7][129] = 16'sd-23;
        fc1_weights[7][130] = 16'sd45;
        fc1_weights[7][131] = 16'sd50;
        fc1_weights[7][132] = 16'sd27;
        fc1_weights[7][133] = 16'sd18;
        fc1_weights[7][134] = 16'sd16;
        fc1_weights[7][135] = 16'sd28;
        fc1_weights[7][136] = 16'sd6;
        fc1_weights[7][137] = 16'sd-6;
        fc1_weights[7][138] = 16'sd-5;
        fc1_weights[7][139] = 16'sd-20;
        fc1_weights[7][140] = 16'sd35;
        fc1_weights[7][141] = 16'sd24;
        fc1_weights[7][142] = 16'sd-14;
        fc1_weights[7][143] = 16'sd-5;
        fc1_weights[7][144] = 16'sd6;
        fc1_weights[7][145] = 16'sd-1;
        fc1_weights[7][146] = 16'sd-12;
        fc1_weights[7][147] = 16'sd-19;
        fc1_weights[7][148] = 16'sd-17;
        fc1_weights[7][149] = 16'sd-28;
        fc1_weights[7][150] = 16'sd-15;
        fc1_weights[7][151] = 16'sd-14;
        fc1_weights[7][152] = 16'sd-14;
        fc1_weights[7][153] = 16'sd-12;
        fc1_weights[7][154] = 16'sd-11;
        fc1_weights[7][155] = 16'sd-5;
        fc1_weights[7][156] = 16'sd-8;
        fc1_weights[7][157] = 16'sd0;
        fc1_weights[7][158] = 16'sd18;
        fc1_weights[7][159] = 16'sd21;
        fc1_weights[7][160] = 16'sd15;
        fc1_weights[7][161] = 16'sd-16;
        fc1_weights[7][162] = 16'sd-23;
        fc1_weights[7][163] = 16'sd-43;
        fc1_weights[7][164] = 16'sd-18;
        fc1_weights[7][165] = 16'sd-1;
        fc1_weights[7][166] = 16'sd0;
        fc1_weights[7][167] = 16'sd-13;
        fc1_weights[7][168] = 16'sd-16;
        fc1_weights[7][169] = 16'sd-8;
        fc1_weights[7][170] = 16'sd-28;
        fc1_weights[7][171] = 16'sd-14;
        fc1_weights[7][172] = 16'sd-13;
        fc1_weights[7][173] = 16'sd-5;
        fc1_weights[7][174] = 16'sd-10;
        fc1_weights[7][175] = 16'sd3;
        fc1_weights[7][176] = 16'sd-6;
        fc1_weights[7][177] = 16'sd13;
        fc1_weights[7][178] = 16'sd-1;
        fc1_weights[7][179] = 16'sd-15;
        fc1_weights[7][180] = 16'sd-18;
        fc1_weights[7][181] = 16'sd5;
        fc1_weights[7][182] = 16'sd11;
        fc1_weights[7][183] = 16'sd12;
        fc1_weights[7][184] = 16'sd10;
        fc1_weights[7][185] = 16'sd-13;
        fc1_weights[7][186] = 16'sd-30;
        fc1_weights[7][187] = 16'sd-23;
        fc1_weights[7][188] = 16'sd3;
        fc1_weights[7][189] = 16'sd-29;
        fc1_weights[7][190] = 16'sd-21;
        fc1_weights[7][191] = 16'sd-15;
        fc1_weights[7][192] = 16'sd2;
        fc1_weights[7][193] = 16'sd5;
        fc1_weights[7][194] = 16'sd-20;
        fc1_weights[7][195] = 16'sd-13;
        fc1_weights[7][196] = 16'sd-17;
        fc1_weights[7][197] = 16'sd-12;
        fc1_weights[7][198] = 16'sd6;
        fc1_weights[7][199] = 16'sd-27;
        fc1_weights[7][200] = 16'sd-22;
        fc1_weights[7][201] = 16'sd-15;
        fc1_weights[7][202] = 16'sd-4;
        fc1_weights[7][203] = 16'sd-9;
        fc1_weights[7][204] = 16'sd6;
        fc1_weights[7][205] = 16'sd0;
        fc1_weights[7][206] = 16'sd5;
        fc1_weights[7][207] = 16'sd6;
        fc1_weights[8][0] = 16'sd-27;
        fc1_weights[8][1] = 16'sd-39;
        fc1_weights[8][2] = 16'sd3;
        fc1_weights[8][3] = 16'sd63;
        fc1_weights[8][4] = 16'sd26;
        fc1_weights[8][5] = 16'sd-10;
        fc1_weights[8][6] = 16'sd-32;
        fc1_weights[8][7] = 16'sd-88;
        fc1_weights[8][8] = 16'sd32;
        fc1_weights[8][9] = 16'sd59;
        fc1_weights[8][10] = 16'sd-57;
        fc1_weights[8][11] = 16'sd64;
        fc1_weights[8][12] = 16'sd119;
        fc1_weights[8][13] = 16'sd51;
        fc1_weights[8][14] = 16'sd10;
        fc1_weights[8][15] = 16'sd-76;
        fc1_weights[8][16] = 16'sd-30;
        fc1_weights[8][17] = 16'sd-41;
        fc1_weights[8][18] = 16'sd-14;
        fc1_weights[8][19] = 16'sd7;
        fc1_weights[8][20] = 16'sd-30;
        fc1_weights[8][21] = 16'sd22;
        fc1_weights[8][22] = 16'sd31;
        fc1_weights[8][23] = 16'sd71;
        fc1_weights[8][24] = 16'sd-18;
        fc1_weights[8][25] = 16'sd-49;
        fc1_weights[8][26] = 16'sd5;
        fc1_weights[8][27] = 16'sd30;
        fc1_weights[8][28] = 16'sd36;
        fc1_weights[8][29] = 16'sd-18;
        fc1_weights[8][30] = 16'sd-47;
        fc1_weights[8][31] = 16'sd-45;
        fc1_weights[8][32] = 16'sd-13;
        fc1_weights[8][33] = 16'sd87;
        fc1_weights[8][34] = 16'sd-24;
        fc1_weights[8][35] = 16'sd-66;
        fc1_weights[8][36] = 16'sd-149;
        fc1_weights[8][37] = 16'sd-149;
        fc1_weights[8][38] = 16'sd-32;
        fc1_weights[8][39] = 16'sd64;
        fc1_weights[8][40] = 16'sd-139;
        fc1_weights[8][41] = 16'sd38;
        fc1_weights[8][42] = 16'sd81;
        fc1_weights[8][43] = 16'sd-60;
        fc1_weights[8][44] = 16'sd-72;
        fc1_weights[8][45] = 16'sd-33;
        fc1_weights[8][46] = 16'sd10;
        fc1_weights[8][47] = 16'sd-63;
        fc1_weights[8][48] = 16'sd-100;
        fc1_weights[8][49] = 16'sd-76;
        fc1_weights[8][50] = 16'sd58;
        fc1_weights[8][51] = 16'sd78;
        fc1_weights[8][52] = 16'sd-19;
        fc1_weights[8][53] = 16'sd-55;
        fc1_weights[8][54] = 16'sd-3;
        fc1_weights[8][55] = 16'sd-68;
        fc1_weights[8][56] = 16'sd-23;
        fc1_weights[8][57] = 16'sd-136;
        fc1_weights[8][58] = 16'sd-11;
        fc1_weights[8][59] = 16'sd18;
        fc1_weights[8][60] = 16'sd-40;
        fc1_weights[8][61] = 16'sd-88;
        fc1_weights[8][62] = 16'sd49;
        fc1_weights[8][63] = 16'sd-59;
        fc1_weights[8][64] = 16'sd17;
        fc1_weights[8][65] = 16'sd38;
        fc1_weights[8][66] = 16'sd-25;
        fc1_weights[8][67] = 16'sd24;
        fc1_weights[8][68] = 16'sd81;
        fc1_weights[8][69] = 16'sd-40;
        fc1_weights[8][70] = 16'sd-54;
        fc1_weights[8][71] = 16'sd-26;
        fc1_weights[8][72] = 16'sd-14;
        fc1_weights[8][73] = 16'sd21;
        fc1_weights[8][74] = 16'sd-34;
        fc1_weights[8][75] = 16'sd3;
        fc1_weights[8][76] = 16'sd-40;
        fc1_weights[8][77] = 16'sd56;
        fc1_weights[8][78] = 16'sd-113;
        fc1_weights[8][79] = 16'sd-110;
        fc1_weights[8][80] = 16'sd-11;
        fc1_weights[8][81] = 16'sd-36;
        fc1_weights[8][82] = 16'sd57;
        fc1_weights[8][83] = 16'sd13;
        fc1_weights[8][84] = 16'sd49;
        fc1_weights[8][85] = 16'sd62;
        fc1_weights[8][86] = 16'sd93;
        fc1_weights[8][87] = 16'sd-35;
        fc1_weights[8][88] = 16'sd12;
        fc1_weights[8][89] = 16'sd-62;
        fc1_weights[8][90] = 16'sd-31;
        fc1_weights[8][91] = 16'sd-17;
        fc1_weights[8][92] = 16'sd-32;
        fc1_weights[8][93] = 16'sd-20;
        fc1_weights[8][94] = 16'sd24;
        fc1_weights[8][95] = 16'sd36;
        fc1_weights[8][96] = 16'sd21;
        fc1_weights[8][97] = 16'sd5;
        fc1_weights[8][98] = 16'sd12;
        fc1_weights[8][99] = 16'sd-61;
        fc1_weights[8][100] = 16'sd-50;
        fc1_weights[8][101] = 16'sd-71;
        fc1_weights[8][102] = 16'sd16;
        fc1_weights[8][103] = 16'sd29;
        fc1_weights[8][104] = 16'sd-61;
        fc1_weights[8][105] = 16'sd-16;
        fc1_weights[8][106] = 16'sd15;
        fc1_weights[8][107] = 16'sd-112;
        fc1_weights[8][108] = 16'sd-128;
        fc1_weights[8][109] = 16'sd-53;
        fc1_weights[8][110] = 16'sd1;
        fc1_weights[8][111] = 16'sd1;
        fc1_weights[8][112] = 16'sd-87;
        fc1_weights[8][113] = 16'sd-56;
        fc1_weights[8][114] = 16'sd-63;
        fc1_weights[8][115] = 16'sd33;
        fc1_weights[8][116] = 16'sd-11;
        fc1_weights[8][117] = 16'sd-24;
        fc1_weights[8][118] = 16'sd-17;
        fc1_weights[8][119] = 16'sd-16;
        fc1_weights[8][120] = 16'sd41;
        fc1_weights[8][121] = 16'sd9;
        fc1_weights[8][122] = 16'sd1;
        fc1_weights[8][123] = 16'sd-5;
        fc1_weights[8][124] = 16'sd-38;
        fc1_weights[8][125] = 16'sd1;
        fc1_weights[8][126] = 16'sd61;
        fc1_weights[8][127] = 16'sd-73;
        fc1_weights[8][128] = 16'sd-7;
        fc1_weights[8][129] = 16'sd176;
        fc1_weights[8][130] = 16'sd-8;
        fc1_weights[8][131] = 16'sd-31;
        fc1_weights[8][132] = 16'sd-17;
        fc1_weights[8][133] = 16'sd-44;
        fc1_weights[8][134] = 16'sd-9;
        fc1_weights[8][135] = 16'sd-16;
        fc1_weights[8][136] = 16'sd-49;
        fc1_weights[8][137] = 16'sd-19;
        fc1_weights[8][138] = 16'sd-80;
        fc1_weights[8][139] = 16'sd7;
        fc1_weights[8][140] = 16'sd-19;
        fc1_weights[8][141] = 16'sd97;
        fc1_weights[8][142] = 16'sd-55;
        fc1_weights[8][143] = 16'sd-45;
        fc1_weights[8][144] = 16'sd-74;
        fc1_weights[8][145] = 16'sd31;
        fc1_weights[8][146] = 16'sd-10;
        fc1_weights[8][147] = 16'sd-91;
        fc1_weights[8][148] = 16'sd-76;
        fc1_weights[8][149] = 16'sd-17;
        fc1_weights[8][150] = 16'sd-15;
        fc1_weights[8][151] = 16'sd6;
        fc1_weights[8][152] = 16'sd-49;
        fc1_weights[8][153] = 16'sd-56;
        fc1_weights[8][154] = 16'sd29;
        fc1_weights[8][155] = 16'sd-69;
        fc1_weights[8][156] = 16'sd18;
        fc1_weights[8][157] = 16'sd-4;
        fc1_weights[8][158] = 16'sd-51;
        fc1_weights[8][159] = 16'sd10;
        fc1_weights[8][160] = 16'sd91;
        fc1_weights[8][161] = 16'sd106;
        fc1_weights[8][162] = 16'sd-33;
        fc1_weights[8][163] = 16'sd58;
        fc1_weights[8][164] = 16'sd-57;
        fc1_weights[8][165] = 16'sd-19;
        fc1_weights[8][166] = 16'sd-105;
        fc1_weights[8][167] = 16'sd-67;
        fc1_weights[8][168] = 16'sd-68;
        fc1_weights[8][169] = 16'sd-7;
        fc1_weights[8][170] = 16'sd-9;
        fc1_weights[8][171] = 16'sd5;
        fc1_weights[8][172] = 16'sd-19;
        fc1_weights[8][173] = 16'sd88;
        fc1_weights[8][174] = 16'sd103;
        fc1_weights[8][175] = 16'sd9;
        fc1_weights[8][176] = 16'sd18;
        fc1_weights[8][177] = 16'sd-40;
        fc1_weights[8][178] = 16'sd-9;
        fc1_weights[8][179] = 16'sd-35;
        fc1_weights[8][180] = 16'sd-17;
        fc1_weights[8][181] = 16'sd-67;
        fc1_weights[8][182] = 16'sd-8;
        fc1_weights[8][183] = 16'sd-27;
        fc1_weights[8][184] = 16'sd57;
        fc1_weights[8][185] = 16'sd-25;
        fc1_weights[8][186] = 16'sd-23;
        fc1_weights[8][187] = 16'sd-11;
        fc1_weights[8][188] = 16'sd55;
        fc1_weights[8][189] = 16'sd7;
        fc1_weights[8][190] = 16'sd-50;
        fc1_weights[8][191] = 16'sd-81;
        fc1_weights[8][192] = 16'sd11;
        fc1_weights[8][193] = 16'sd-40;
        fc1_weights[8][194] = 16'sd-55;
        fc1_weights[8][195] = 16'sd4;
        fc1_weights[8][196] = 16'sd48;
        fc1_weights[8][197] = 16'sd-100;
        fc1_weights[8][198] = 16'sd46;
        fc1_weights[8][199] = 16'sd-11;
        fc1_weights[8][200] = 16'sd28;
        fc1_weights[8][201] = 16'sd6;
        fc1_weights[8][202] = 16'sd8;
        fc1_weights[8][203] = 16'sd-12;
        fc1_weights[8][204] = 16'sd-47;
        fc1_weights[8][205] = 16'sd-55;
        fc1_weights[8][206] = 16'sd82;
        fc1_weights[8][207] = 16'sd-26;
        fc1_weights[9][0] = 16'sd5;
        fc1_weights[9][1] = 16'sd8;
        fc1_weights[9][2] = 16'sd15;
        fc1_weights[9][3] = 16'sd1;
        fc1_weights[9][4] = 16'sd7;
        fc1_weights[9][5] = 16'sd-21;
        fc1_weights[9][6] = 16'sd-1;
        fc1_weights[9][7] = 16'sd-20;
        fc1_weights[9][8] = 16'sd-32;
        fc1_weights[9][9] = 16'sd4;
        fc1_weights[9][10] = 16'sd-23;
        fc1_weights[9][11] = 16'sd19;
        fc1_weights[9][12] = 16'sd-16;
        fc1_weights[9][13] = 16'sd-9;
        fc1_weights[9][14] = 16'sd9;
        fc1_weights[9][15] = 16'sd-15;
        fc1_weights[9][16] = 16'sd29;
        fc1_weights[9][17] = 16'sd53;
        fc1_weights[9][18] = 16'sd8;
        fc1_weights[9][19] = 16'sd50;
        fc1_weights[9][20] = 16'sd52;
        fc1_weights[9][21] = 16'sd9;
        fc1_weights[9][22] = 16'sd11;
        fc1_weights[9][23] = 16'sd30;
        fc1_weights[9][24] = 16'sd12;
        fc1_weights[9][25] = 16'sd-8;
        fc1_weights[9][26] = 16'sd22;
        fc1_weights[9][27] = 16'sd2;
        fc1_weights[9][28] = 16'sd23;
        fc1_weights[9][29] = 16'sd32;
        fc1_weights[9][30] = 16'sd-25;
        fc1_weights[9][31] = 16'sd-23;
        fc1_weights[9][32] = 16'sd-7;
        fc1_weights[9][33] = 16'sd48;
        fc1_weights[9][34] = 16'sd1;
        fc1_weights[9][35] = 16'sd-3;
        fc1_weights[9][36] = 16'sd-3;
        fc1_weights[9][37] = 16'sd-32;
        fc1_weights[9][38] = 16'sd-15;
        fc1_weights[9][39] = 16'sd-27;
        fc1_weights[9][40] = 16'sd36;
        fc1_weights[9][41] = 16'sd-6;
        fc1_weights[9][42] = 16'sd17;
        fc1_weights[9][43] = 16'sd58;
        fc1_weights[9][44] = 16'sd44;
        fc1_weights[9][45] = 16'sd64;
        fc1_weights[9][46] = 16'sd39;
        fc1_weights[9][47] = 16'sd4;
        fc1_weights[9][48] = 16'sd8;
        fc1_weights[9][49] = 16'sd-18;
        fc1_weights[9][50] = 16'sd4;
        fc1_weights[9][51] = 16'sd-28;
        fc1_weights[9][52] = 16'sd13;
        fc1_weights[9][53] = 16'sd-13;
        fc1_weights[9][54] = 16'sd18;
        fc1_weights[9][55] = 16'sd30;
        fc1_weights[9][56] = 16'sd4;
        fc1_weights[9][57] = 16'sd29;
        fc1_weights[9][58] = 16'sd33;
        fc1_weights[9][59] = 16'sd38;
        fc1_weights[9][60] = 16'sd4;
        fc1_weights[9][61] = 16'sd-20;
        fc1_weights[9][62] = 16'sd-10;
        fc1_weights[9][63] = 16'sd1;
        fc1_weights[9][64] = 16'sd-16;
        fc1_weights[9][65] = 16'sd-27;
        fc1_weights[9][66] = 16'sd-29;
        fc1_weights[9][67] = 16'sd-34;
        fc1_weights[9][68] = 16'sd-4;
        fc1_weights[9][69] = 16'sd10;
        fc1_weights[9][70] = 16'sd-11;
        fc1_weights[9][71] = 16'sd25;
        fc1_weights[9][72] = 16'sd1;
        fc1_weights[9][73] = 16'sd-14;
        fc1_weights[9][74] = 16'sd-10;
        fc1_weights[9][75] = 16'sd-27;
        fc1_weights[9][76] = 16'sd-4;
        fc1_weights[9][77] = 16'sd-11;
        fc1_weights[9][78] = 16'sd9;
        fc1_weights[9][79] = 16'sd23;
        fc1_weights[9][80] = 16'sd8;
        fc1_weights[9][81] = 16'sd9;
        fc1_weights[9][82] = 16'sd35;
        fc1_weights[9][83] = 16'sd-2;
        fc1_weights[9][84] = 16'sd47;
        fc1_weights[9][85] = 16'sd9;
        fc1_weights[9][86] = 16'sd-7;
        fc1_weights[9][87] = 16'sd-16;
        fc1_weights[9][88] = 16'sd-14;
        fc1_weights[9][89] = 16'sd-29;
        fc1_weights[9][90] = 16'sd-48;
        fc1_weights[9][91] = 16'sd-40;
        fc1_weights[9][92] = 16'sd-30;
        fc1_weights[9][93] = 16'sd-7;
        fc1_weights[9][94] = 16'sd8;
        fc1_weights[9][95] = 16'sd6;
        fc1_weights[9][96] = 16'sd-17;
        fc1_weights[9][97] = 16'sd7;
        fc1_weights[9][98] = 16'sd-4;
        fc1_weights[9][99] = 16'sd-39;
        fc1_weights[9][100] = 16'sd-19;
        fc1_weights[9][101] = 16'sd-14;
        fc1_weights[9][102] = 16'sd-20;
        fc1_weights[9][103] = 16'sd12;
        fc1_weights[9][104] = 16'sd12;
        fc1_weights[9][105] = 16'sd5;
        fc1_weights[9][106] = 16'sd-21;
        fc1_weights[9][107] = 16'sd-10;
        fc1_weights[9][108] = 16'sd-10;
        fc1_weights[9][109] = 16'sd-6;
        fc1_weights[9][110] = 16'sd-4;
        fc1_weights[9][111] = 16'sd22;
        fc1_weights[9][112] = 16'sd-57;
        fc1_weights[9][113] = 16'sd-26;
        fc1_weights[9][114] = 16'sd12;
        fc1_weights[9][115] = 16'sd0;
        fc1_weights[9][116] = 16'sd64;
        fc1_weights[9][117] = 16'sd-56;
        fc1_weights[9][118] = 16'sd-41;
        fc1_weights[9][119] = 16'sd-33;
        fc1_weights[9][120] = 16'sd-19;
        fc1_weights[9][121] = 16'sd-18;
        fc1_weights[9][122] = 16'sd-15;
        fc1_weights[9][123] = 16'sd9;
        fc1_weights[9][124] = 16'sd20;
        fc1_weights[9][125] = 16'sd23;
        fc1_weights[9][126] = 16'sd5;
        fc1_weights[9][127] = 16'sd-43;
        fc1_weights[9][128] = 16'sd-21;
        fc1_weights[9][129] = 16'sd-10;
        fc1_weights[9][130] = 16'sd15;
        fc1_weights[9][131] = 16'sd-41;
        fc1_weights[9][132] = 16'sd-45;
        fc1_weights[9][133] = 16'sd-56;
        fc1_weights[9][134] = 16'sd-29;
        fc1_weights[9][135] = 16'sd-21;
        fc1_weights[9][136] = 16'sd-18;
        fc1_weights[9][137] = 16'sd-9;
        fc1_weights[9][138] = 16'sd15;
        fc1_weights[9][139] = 16'sd62;
        fc1_weights[9][140] = 16'sd38;
        fc1_weights[9][141] = 16'sd3;
        fc1_weights[9][142] = 16'sd-5;
        fc1_weights[9][143] = 16'sd28;
        fc1_weights[9][144] = 16'sd-10;
        fc1_weights[9][145] = 16'sd11;
        fc1_weights[9][146] = 16'sd16;
        fc1_weights[9][147] = 16'sd-6;
        fc1_weights[9][148] = 16'sd0;
        fc1_weights[9][149] = 16'sd-8;
        fc1_weights[9][150] = 16'sd2;
        fc1_weights[9][151] = 16'sd-6;
        fc1_weights[9][152] = 16'sd-20;
        fc1_weights[9][153] = 16'sd-3;
        fc1_weights[9][154] = 16'sd6;
        fc1_weights[9][155] = 16'sd0;
        fc1_weights[9][156] = 16'sd7;
        fc1_weights[9][157] = 16'sd-21;
        fc1_weights[9][158] = 16'sd8;
        fc1_weights[9][159] = 16'sd13;
        fc1_weights[9][160] = 16'sd-9;
        fc1_weights[9][161] = 16'sd-12;
        fc1_weights[9][162] = 16'sd-48;
        fc1_weights[9][163] = 16'sd-31;
        fc1_weights[9][164] = 16'sd38;
        fc1_weights[9][165] = 16'sd28;
        fc1_weights[9][166] = 16'sd33;
        fc1_weights[9][167] = 16'sd1;
        fc1_weights[9][168] = 16'sd-14;
        fc1_weights[9][169] = 16'sd-26;
        fc1_weights[9][170] = 16'sd-49;
        fc1_weights[9][171] = 16'sd-2;
        fc1_weights[9][172] = 16'sd-19;
        fc1_weights[9][173] = 16'sd-13;
        fc1_weights[9][174] = 16'sd-21;
        fc1_weights[9][175] = 16'sd-27;
        fc1_weights[9][176] = 16'sd4;
        fc1_weights[9][177] = 16'sd2;
        fc1_weights[9][178] = 16'sd-5;
        fc1_weights[9][179] = 16'sd13;
        fc1_weights[9][180] = 16'sd-1;
        fc1_weights[9][181] = 16'sd-22;
        fc1_weights[9][182] = 16'sd1;
        fc1_weights[9][183] = 16'sd-21;
        fc1_weights[9][184] = 16'sd-6;
        fc1_weights[9][185] = 16'sd-50;
        fc1_weights[9][186] = 16'sd-22;
        fc1_weights[9][187] = 16'sd-16;
        fc1_weights[9][188] = 16'sd44;
        fc1_weights[9][189] = 16'sd-7;
        fc1_weights[9][190] = 16'sd-2;
        fc1_weights[9][191] = 16'sd-1;
        fc1_weights[9][192] = 16'sd-7;
        fc1_weights[9][193] = 16'sd-1;
        fc1_weights[9][194] = 16'sd-6;
        fc1_weights[9][195] = 16'sd-32;
        fc1_weights[9][196] = 16'sd-18;
        fc1_weights[9][197] = 16'sd-40;
        fc1_weights[9][198] = 16'sd8;
        fc1_weights[9][199] = 16'sd-12;
        fc1_weights[9][200] = 16'sd-12;
        fc1_weights[9][201] = 16'sd2;
        fc1_weights[9][202] = 16'sd-12;
        fc1_weights[9][203] = 16'sd-13;
        fc1_weights[9][204] = 16'sd9;
        fc1_weights[9][205] = 16'sd12;
        fc1_weights[9][206] = 16'sd-5;
        fc1_weights[9][207] = 16'sd-2;
        fc1_weights[10][0] = 16'sd-31;
        fc1_weights[10][1] = 16'sd-23;
        fc1_weights[10][2] = 16'sd-15;
        fc1_weights[10][3] = 16'sd12;
        fc1_weights[10][4] = 16'sd10;
        fc1_weights[10][5] = 16'sd17;
        fc1_weights[10][6] = 16'sd1;
        fc1_weights[10][7] = 16'sd5;
        fc1_weights[10][8] = 16'sd32;
        fc1_weights[10][9] = 16'sd5;
        fc1_weights[10][10] = 16'sd14;
        fc1_weights[10][11] = 16'sd5;
        fc1_weights[10][12] = 16'sd-1;
        fc1_weights[10][13] = 16'sd-14;
        fc1_weights[10][14] = 16'sd-56;
        fc1_weights[10][15] = 16'sd17;
        fc1_weights[10][16] = 16'sd-11;
        fc1_weights[10][17] = 16'sd14;
        fc1_weights[10][18] = 16'sd6;
        fc1_weights[10][19] = 16'sd26;
        fc1_weights[10][20] = 16'sd9;
        fc1_weights[10][21] = 16'sd3;
        fc1_weights[10][22] = 16'sd7;
        fc1_weights[10][23] = 16'sd-9;
        fc1_weights[10][24] = 16'sd15;
        fc1_weights[10][25] = 16'sd20;
        fc1_weights[10][26] = 16'sd-9;
        fc1_weights[10][27] = 16'sd-12;
        fc1_weights[10][28] = 16'sd-37;
        fc1_weights[10][29] = 16'sd-8;
        fc1_weights[10][30] = 16'sd24;
        fc1_weights[10][31] = 16'sd14;
        fc1_weights[10][32] = 16'sd24;
        fc1_weights[10][33] = 16'sd-30;
        fc1_weights[10][34] = 16'sd5;
        fc1_weights[10][35] = 16'sd-14;
        fc1_weights[10][36] = 16'sd27;
        fc1_weights[10][37] = 16'sd9;
        fc1_weights[10][38] = 16'sd27;
        fc1_weights[10][39] = 16'sd33;
        fc1_weights[10][40] = 16'sd3;
        fc1_weights[10][41] = 16'sd4;
        fc1_weights[10][42] = 16'sd19;
        fc1_weights[10][43] = 16'sd15;
        fc1_weights[10][44] = 16'sd54;
        fc1_weights[10][45] = 16'sd18;
        fc1_weights[10][46] = 16'sd16;
        fc1_weights[10][47] = 16'sd-12;
        fc1_weights[10][48] = 16'sd-1;
        fc1_weights[10][49] = 16'sd27;
        fc1_weights[10][50] = 16'sd-3;
        fc1_weights[10][51] = 16'sd-4;
        fc1_weights[10][52] = 16'sd-31;
        fc1_weights[10][53] = 16'sd-22;
        fc1_weights[10][54] = 16'sd-11;
        fc1_weights[10][55] = 16'sd-14;
        fc1_weights[10][56] = 16'sd-19;
        fc1_weights[10][57] = 16'sd-2;
        fc1_weights[10][58] = 16'sd-15;
        fc1_weights[10][59] = 16'sd14;
        fc1_weights[10][60] = 16'sd40;
        fc1_weights[10][61] = 16'sd31;
        fc1_weights[10][62] = 16'sd17;
        fc1_weights[10][63] = 16'sd26;
        fc1_weights[10][64] = 16'sd65;
        fc1_weights[10][65] = 16'sd22;
        fc1_weights[10][66] = 16'sd22;
        fc1_weights[10][67] = 16'sd-10;
        fc1_weights[10][68] = 16'sd9;
        fc1_weights[10][69] = 16'sd-13;
        fc1_weights[10][70] = 16'sd32;
        fc1_weights[10][71] = 16'sd18;
        fc1_weights[10][72] = 16'sd-9;
        fc1_weights[10][73] = 16'sd14;
        fc1_weights[10][74] = 16'sd-6;
        fc1_weights[10][75] = 16'sd20;
        fc1_weights[10][76] = 16'sd11;
        fc1_weights[10][77] = 16'sd1;
        fc1_weights[10][78] = 16'sd-2;
        fc1_weights[10][79] = 16'sd18;
        fc1_weights[10][80] = 16'sd41;
        fc1_weights[10][81] = 16'sd0;
        fc1_weights[10][82] = 16'sd-6;
        fc1_weights[10][83] = 16'sd-5;
        fc1_weights[10][84] = 16'sd-38;
        fc1_weights[10][85] = 16'sd-5;
        fc1_weights[10][86] = 16'sd-14;
        fc1_weights[10][87] = 16'sd44;
        fc1_weights[10][88] = 16'sd31;
        fc1_weights[10][89] = 16'sd37;
        fc1_weights[10][90] = 16'sd68;
        fc1_weights[10][91] = 16'sd41;
        fc1_weights[10][92] = 16'sd5;
        fc1_weights[10][93] = 16'sd-8;
        fc1_weights[10][94] = 16'sd-6;
        fc1_weights[10][95] = 16'sd-6;
        fc1_weights[10][96] = 16'sd0;
        fc1_weights[10][97] = 16'sd8;
        fc1_weights[10][98] = 16'sd-13;
        fc1_weights[10][99] = 16'sd1;
        fc1_weights[10][100] = 16'sd-12;
        fc1_weights[10][101] = 16'sd-21;
        fc1_weights[10][102] = 16'sd-22;
        fc1_weights[10][103] = 16'sd0;
        fc1_weights[10][104] = 16'sd-9;
        fc1_weights[10][105] = 16'sd3;
        fc1_weights[10][106] = 16'sd17;
        fc1_weights[10][107] = 16'sd6;
        fc1_weights[10][108] = 16'sd20;
        fc1_weights[10][109] = 16'sd45;
        fc1_weights[10][110] = 16'sd25;
        fc1_weights[10][111] = 16'sd26;
        fc1_weights[10][112] = 16'sd36;
        fc1_weights[10][113] = 16'sd24;
        fc1_weights[10][114] = 16'sd2;
        fc1_weights[10][115] = 16'sd-8;
        fc1_weights[10][116] = 16'sd-7;
        fc1_weights[10][117] = 16'sd60;
        fc1_weights[10][118] = 16'sd40;
        fc1_weights[10][119] = 16'sd8;
        fc1_weights[10][120] = 16'sd-3;
        fc1_weights[10][121] = 16'sd14;
        fc1_weights[10][122] = 16'sd34;
        fc1_weights[10][123] = 16'sd42;
        fc1_weights[10][124] = 16'sd-5;
        fc1_weights[10][125] = 16'sd10;
        fc1_weights[10][126] = 16'sd-4;
        fc1_weights[10][127] = 16'sd14;
        fc1_weights[10][128] = 16'sd17;
        fc1_weights[10][129] = 16'sd28;
        fc1_weights[10][130] = 16'sd4;
        fc1_weights[10][131] = 16'sd37;
        fc1_weights[10][132] = 16'sd25;
        fc1_weights[10][133] = 16'sd32;
        fc1_weights[10][134] = 16'sd27;
        fc1_weights[10][135] = 16'sd57;
        fc1_weights[10][136] = 16'sd34;
        fc1_weights[10][137] = 16'sd32;
        fc1_weights[10][138] = 16'sd17;
        fc1_weights[10][139] = 16'sd4;
        fc1_weights[10][140] = 16'sd-12;
        fc1_weights[10][141] = 16'sd-11;
        fc1_weights[10][142] = 16'sd13;
        fc1_weights[10][143] = 16'sd14;
        fc1_weights[10][144] = 16'sd8;
        fc1_weights[10][145] = 16'sd-6;
        fc1_weights[10][146] = 16'sd-18;
        fc1_weights[10][147] = 16'sd-18;
        fc1_weights[10][148] = 16'sd-18;
        fc1_weights[10][149] = 16'sd-11;
        fc1_weights[10][150] = 16'sd0;
        fc1_weights[10][151] = 16'sd24;
        fc1_weights[10][152] = 16'sd-13;
        fc1_weights[10][153] = 16'sd6;
        fc1_weights[10][154] = 16'sd0;
        fc1_weights[10][155] = 16'sd-11;
        fc1_weights[10][156] = 16'sd26;
        fc1_weights[10][157] = 16'sd34;
        fc1_weights[10][158] = 16'sd-7;
        fc1_weights[10][159] = 16'sd10;
        fc1_weights[10][160] = 16'sd-25;
        fc1_weights[10][161] = 16'sd-9;
        fc1_weights[10][162] = 16'sd12;
        fc1_weights[10][163] = 16'sd-3;
        fc1_weights[10][164] = 16'sd-18;
        fc1_weights[10][165] = 16'sd-47;
        fc1_weights[10][166] = 16'sd-29;
        fc1_weights[10][167] = 16'sd-13;
        fc1_weights[10][168] = 16'sd-5;
        fc1_weights[10][169] = 16'sd29;
        fc1_weights[10][170] = 16'sd49;
        fc1_weights[10][171] = 16'sd0;
        fc1_weights[10][172] = 16'sd-6;
        fc1_weights[10][173] = 16'sd-23;
        fc1_weights[10][174] = 16'sd-25;
        fc1_weights[10][175] = 16'sd-9;
        fc1_weights[10][176] = 16'sd-22;
        fc1_weights[10][177] = 16'sd-8;
        fc1_weights[10][178] = 16'sd-8;
        fc1_weights[10][179] = 16'sd9;
        fc1_weights[10][180] = 16'sd1;
        fc1_weights[10][181] = 16'sd-7;
        fc1_weights[10][182] = 16'sd2;
        fc1_weights[10][183] = 16'sd13;
        fc1_weights[10][184] = 16'sd14;
        fc1_weights[10][185] = 16'sd-6;
        fc1_weights[10][186] = 16'sd-17;
        fc1_weights[10][187] = 16'sd-5;
        fc1_weights[10][188] = 16'sd-18;
        fc1_weights[10][189] = 16'sd10;
        fc1_weights[10][190] = 16'sd-5;
        fc1_weights[10][191] = 16'sd-25;
        fc1_weights[10][192] = 16'sd-29;
        fc1_weights[10][193] = 16'sd-19;
        fc1_weights[10][194] = 16'sd-17;
        fc1_weights[10][195] = 16'sd-13;
        fc1_weights[10][196] = 16'sd8;
        fc1_weights[10][197] = 16'sd40;
        fc1_weights[10][198] = 16'sd-23;
        fc1_weights[10][199] = 16'sd-14;
        fc1_weights[10][200] = 16'sd-7;
        fc1_weights[10][201] = 16'sd2;
        fc1_weights[10][202] = 16'sd12;
        fc1_weights[10][203] = 16'sd-7;
        fc1_weights[10][204] = 16'sd9;
        fc1_weights[10][205] = 16'sd-21;
        fc1_weights[10][206] = 16'sd-25;
        fc1_weights[10][207] = 16'sd-18;
        fc1_weights[11][0] = 16'sd-10;
        fc1_weights[11][1] = 16'sd25;
        fc1_weights[11][2] = 16'sd-31;
        fc1_weights[11][3] = 16'sd0;
        fc1_weights[11][4] = 16'sd44;
        fc1_weights[11][5] = 16'sd13;
        fc1_weights[11][6] = 16'sd8;
        fc1_weights[11][7] = 16'sd56;
        fc1_weights[11][8] = 16'sd27;
        fc1_weights[11][9] = 16'sd10;
        fc1_weights[11][10] = 16'sd7;
        fc1_weights[11][11] = 16'sd5;
        fc1_weights[11][12] = 16'sd90;
        fc1_weights[11][13] = 16'sd69;
        fc1_weights[11][14] = 16'sd33;
        fc1_weights[11][15] = 16'sd28;
        fc1_weights[11][16] = 16'sd13;
        fc1_weights[11][17] = 16'sd8;
        fc1_weights[11][18] = 16'sd22;
        fc1_weights[11][19] = 16'sd22;
        fc1_weights[11][20] = 16'sd41;
        fc1_weights[11][21] = 16'sd20;
        fc1_weights[11][22] = 16'sd43;
        fc1_weights[11][23] = 16'sd14;
        fc1_weights[11][24] = 16'sd38;
        fc1_weights[11][25] = 16'sd19;
        fc1_weights[11][26] = 16'sd-2;
        fc1_weights[11][27] = 16'sd-27;
        fc1_weights[11][28] = 16'sd3;
        fc1_weights[11][29] = 16'sd39;
        fc1_weights[11][30] = 16'sd9;
        fc1_weights[11][31] = 16'sd30;
        fc1_weights[11][32] = 16'sd-13;
        fc1_weights[11][33] = 16'sd36;
        fc1_weights[11][34] = 16'sd24;
        fc1_weights[11][35] = 16'sd3;
        fc1_weights[11][36] = 16'sd29;
        fc1_weights[11][37] = 16'sd15;
        fc1_weights[11][38] = 16'sd-6;
        fc1_weights[11][39] = 16'sd84;
        fc1_weights[11][40] = 16'sd5;
        fc1_weights[11][41] = 16'sd17;
        fc1_weights[11][42] = 16'sd3;
        fc1_weights[11][43] = 16'sd37;
        fc1_weights[11][44] = 16'sd-1;
        fc1_weights[11][45] = 16'sd-17;
        fc1_weights[11][46] = 16'sd-23;
        fc1_weights[11][47] = 16'sd29;
        fc1_weights[11][48] = 16'sd-17;
        fc1_weights[11][49] = 16'sd-18;
        fc1_weights[11][50] = 16'sd-18;
        fc1_weights[11][51] = 16'sd1;
        fc1_weights[11][52] = 16'sd43;
        fc1_weights[11][53] = 16'sd-47;
        fc1_weights[11][54] = 16'sd-51;
        fc1_weights[11][55] = 16'sd-29;
        fc1_weights[11][56] = 16'sd-7;
        fc1_weights[11][57] = 16'sd24;
        fc1_weights[11][58] = 16'sd41;
        fc1_weights[11][59] = 16'sd46;
        fc1_weights[11][60] = 16'sd20;
        fc1_weights[11][61] = 16'sd42;
        fc1_weights[11][62] = 16'sd29;
        fc1_weights[11][63] = 16'sd-3;
        fc1_weights[11][64] = 16'sd12;
        fc1_weights[11][65] = 16'sd64;
        fc1_weights[11][66] = 16'sd57;
        fc1_weights[11][67] = 16'sd-16;
        fc1_weights[11][68] = 16'sd-58;
        fc1_weights[11][69] = 16'sd-4;
        fc1_weights[11][70] = 16'sd-24;
        fc1_weights[11][71] = 16'sd1;
        fc1_weights[11][72] = 16'sd24;
        fc1_weights[11][73] = 16'sd7;
        fc1_weights[11][74] = 16'sd30;
        fc1_weights[11][75] = 16'sd8;
        fc1_weights[11][76] = 16'sd-28;
        fc1_weights[11][77] = 16'sd-9;
        fc1_weights[11][78] = 16'sd-7;
        fc1_weights[11][79] = 16'sd-10;
        fc1_weights[11][80] = 16'sd-47;
        fc1_weights[11][81] = 16'sd19;
        fc1_weights[11][82] = 16'sd-8;
        fc1_weights[11][83] = 16'sd59;
        fc1_weights[11][84] = 16'sd2;
        fc1_weights[11][85] = 16'sd14;
        fc1_weights[11][86] = 16'sd8;
        fc1_weights[11][87] = 16'sd41;
        fc1_weights[11][88] = 16'sd36;
        fc1_weights[11][89] = 16'sd-38;
        fc1_weights[11][90] = 16'sd3;
        fc1_weights[11][91] = 16'sd-31;
        fc1_weights[11][92] = 16'sd-30;
        fc1_weights[11][93] = 16'sd-42;
        fc1_weights[11][94] = 16'sd-81;
        fc1_weights[11][95] = 16'sd-19;
        fc1_weights[11][96] = 16'sd-48;
        fc1_weights[11][97] = 16'sd-59;
        fc1_weights[11][98] = 16'sd-14;
        fc1_weights[11][99] = 16'sd-31;
        fc1_weights[11][100] = 16'sd32;
        fc1_weights[11][101] = 16'sd-13;
        fc1_weights[11][102] = 16'sd-16;
        fc1_weights[11][103] = 16'sd-12;
        fc1_weights[11][104] = 16'sd24;
        fc1_weights[11][105] = 16'sd-42;
        fc1_weights[11][106] = 16'sd-18;
        fc1_weights[11][107] = 16'sd4;
        fc1_weights[11][108] = 16'sd-2;
        fc1_weights[11][109] = 16'sd29;
        fc1_weights[11][110] = 16'sd-3;
        fc1_weights[11][111] = 16'sd38;
        fc1_weights[11][112] = 16'sd48;
        fc1_weights[11][113] = 16'sd1;
        fc1_weights[11][114] = 16'sd33;
        fc1_weights[11][115] = 16'sd11;
        fc1_weights[11][116] = 16'sd16;
        fc1_weights[11][117] = 16'sd8;
        fc1_weights[11][118] = 16'sd6;
        fc1_weights[11][119] = 16'sd-25;
        fc1_weights[11][120] = 16'sd-16;
        fc1_weights[11][121] = 16'sd-12;
        fc1_weights[11][122] = 16'sd-14;
        fc1_weights[11][123] = 16'sd-42;
        fc1_weights[11][124] = 16'sd-9;
        fc1_weights[11][125] = 16'sd21;
        fc1_weights[11][126] = 16'sd-10;
        fc1_weights[11][127] = 16'sd-24;
        fc1_weights[11][128] = 16'sd5;
        fc1_weights[11][129] = 16'sd-9;
        fc1_weights[11][130] = 16'sd21;
        fc1_weights[11][131] = 16'sd24;
        fc1_weights[11][132] = 16'sd24;
        fc1_weights[11][133] = 16'sd-17;
        fc1_weights[11][134] = 16'sd-5;
        fc1_weights[11][135] = 16'sd-6;
        fc1_weights[11][136] = 16'sd36;
        fc1_weights[11][137] = 16'sd50;
        fc1_weights[11][138] = 16'sd3;
        fc1_weights[11][139] = 16'sd-42;
        fc1_weights[11][140] = 16'sd21;
        fc1_weights[11][141] = 16'sd63;
        fc1_weights[11][142] = 16'sd-1;
        fc1_weights[11][143] = 16'sd10;
        fc1_weights[11][144] = 16'sd69;
        fc1_weights[11][145] = 16'sd90;
        fc1_weights[11][146] = 16'sd71;
        fc1_weights[11][147] = 16'sd47;
        fc1_weights[11][148] = 16'sd29;
        fc1_weights[11][149] = 16'sd28;
        fc1_weights[11][150] = 16'sd23;
        fc1_weights[11][151] = 16'sd4;
        fc1_weights[11][152] = 16'sd-39;
        fc1_weights[11][153] = 16'sd-21;
        fc1_weights[11][154] = 16'sd9;
        fc1_weights[11][155] = 16'sd-24;
        fc1_weights[11][156] = 16'sd-6;
        fc1_weights[11][157] = 16'sd9;
        fc1_weights[11][158] = 16'sd2;
        fc1_weights[11][159] = 16'sd60;
        fc1_weights[11][160] = 16'sd42;
        fc1_weights[11][161] = 16'sd18;
        fc1_weights[11][162] = 16'sd-19;
        fc1_weights[11][163] = 16'sd1;
        fc1_weights[11][164] = 16'sd-40;
        fc1_weights[11][165] = 16'sd-22;
        fc1_weights[11][166] = 16'sd-6;
        fc1_weights[11][167] = 16'sd20;
        fc1_weights[11][168] = 16'sd-16;
        fc1_weights[11][169] = 16'sd5;
        fc1_weights[11][170] = 16'sd20;
        fc1_weights[11][171] = 16'sd13;
        fc1_weights[11][172] = 16'sd30;
        fc1_weights[11][173] = 16'sd28;
        fc1_weights[11][174] = 16'sd60;
        fc1_weights[11][175] = 16'sd48;
        fc1_weights[11][176] = 16'sd29;
        fc1_weights[11][177] = 16'sd-32;
        fc1_weights[11][178] = 16'sd27;
        fc1_weights[11][179] = 16'sd-36;
        fc1_weights[11][180] = 16'sd-39;
        fc1_weights[11][181] = 16'sd-27;
        fc1_weights[11][182] = 16'sd-44;
        fc1_weights[11][183] = 16'sd-38;
        fc1_weights[11][184] = 16'sd-48;
        fc1_weights[11][185] = 16'sd-14;
        fc1_weights[11][186] = 16'sd-37;
        fc1_weights[11][187] = 16'sd-35;
        fc1_weights[11][188] = 16'sd-2;
        fc1_weights[11][189] = 16'sd-6;
        fc1_weights[11][190] = 16'sd17;
        fc1_weights[11][191] = 16'sd-18;
        fc1_weights[11][192] = 16'sd28;
        fc1_weights[11][193] = 16'sd10;
        fc1_weights[11][194] = 16'sd-13;
        fc1_weights[11][195] = 16'sd6;
        fc1_weights[11][196] = 16'sd-13;
        fc1_weights[11][197] = 16'sd-18;
        fc1_weights[11][198] = 16'sd-12;
        fc1_weights[11][199] = 16'sd-17;
        fc1_weights[11][200] = 16'sd6;
        fc1_weights[11][201] = 16'sd6;
        fc1_weights[11][202] = 16'sd23;
        fc1_weights[11][203] = 16'sd-20;
        fc1_weights[11][204] = 16'sd-39;
        fc1_weights[11][205] = 16'sd-50;
        fc1_weights[11][206] = 16'sd4;
        fc1_weights[11][207] = 16'sd-8;
        fc1_weights[12][0] = 16'sd19;
        fc1_weights[12][1] = 16'sd25;
        fc1_weights[12][2] = 16'sd19;
        fc1_weights[12][3] = 16'sd125;
        fc1_weights[12][4] = 16'sd-1;
        fc1_weights[12][5] = 16'sd77;
        fc1_weights[12][6] = 16'sd66;
        fc1_weights[12][7] = 16'sd46;
        fc1_weights[12][8] = 16'sd47;
        fc1_weights[12][9] = 16'sd77;
        fc1_weights[12][10] = 16'sd28;
        fc1_weights[12][11] = 16'sd59;
        fc1_weights[12][12] = 16'sd131;
        fc1_weights[12][13] = 16'sd20;
        fc1_weights[12][14] = 16'sd115;
        fc1_weights[12][15] = 16'sd5;
        fc1_weights[12][16] = 16'sd-14;
        fc1_weights[12][17] = 16'sd29;
        fc1_weights[12][18] = 16'sd-34;
        fc1_weights[12][19] = 16'sd34;
        fc1_weights[12][20] = 16'sd-42;
        fc1_weights[12][21] = 16'sd13;
        fc1_weights[12][22] = 16'sd12;
        fc1_weights[12][23] = 16'sd0;
        fc1_weights[12][24] = 16'sd-2;
        fc1_weights[12][25] = 16'sd-60;
        fc1_weights[12][26] = 16'sd45;
        fc1_weights[12][27] = 16'sd40;
        fc1_weights[12][28] = 16'sd52;
        fc1_weights[12][29] = 16'sd-31;
        fc1_weights[12][30] = 16'sd-61;
        fc1_weights[12][31] = 16'sd-117;
        fc1_weights[12][32] = 16'sd-11;
        fc1_weights[12][33] = 16'sd92;
        fc1_weights[12][34] = 16'sd38;
        fc1_weights[12][35] = 16'sd21;
        fc1_weights[12][36] = 16'sd-57;
        fc1_weights[12][37] = 16'sd-46;
        fc1_weights[12][38] = 16'sd39;
        fc1_weights[12][39] = 16'sd47;
        fc1_weights[12][40] = 16'sd46;
        fc1_weights[12][41] = 16'sd41;
        fc1_weights[12][42] = 16'sd23;
        fc1_weights[12][43] = 16'sd-8;
        fc1_weights[12][44] = 16'sd-6;
        fc1_weights[12][45] = 16'sd52;
        fc1_weights[12][46] = 16'sd48;
        fc1_weights[12][47] = 16'sd30;
        fc1_weights[12][48] = 16'sd-35;
        fc1_weights[12][49] = 16'sd-64;
        fc1_weights[12][50] = 16'sd29;
        fc1_weights[12][51] = 16'sd47;
        fc1_weights[12][52] = 16'sd30;
        fc1_weights[12][53] = 16'sd-39;
        fc1_weights[12][54] = 16'sd-3;
        fc1_weights[12][55] = 16'sd56;
        fc1_weights[12][56] = 16'sd-22;
        fc1_weights[12][57] = 16'sd-37;
        fc1_weights[12][58] = 16'sd-40;
        fc1_weights[12][59] = 16'sd-1;
        fc1_weights[12][60] = 16'sd-51;
        fc1_weights[12][61] = 16'sd-18;
        fc1_weights[12][62] = 16'sd-19;
        fc1_weights[12][63] = 16'sd-79;
        fc1_weights[12][64] = 16'sd13;
        fc1_weights[12][65] = 16'sd61;
        fc1_weights[12][66] = 16'sd-72;
        fc1_weights[12][67] = 16'sd-40;
        fc1_weights[12][68] = 16'sd36;
        fc1_weights[12][69] = 16'sd-18;
        fc1_weights[12][70] = 16'sd23;
        fc1_weights[12][71] = 16'sd36;
        fc1_weights[12][72] = 16'sd48;
        fc1_weights[12][73] = 16'sd31;
        fc1_weights[12][74] = 16'sd-55;
        fc1_weights[12][75] = 16'sd-37;
        fc1_weights[12][76] = 16'sd-78;
        fc1_weights[12][77] = 16'sd-41;
        fc1_weights[12][78] = 16'sd-39;
        fc1_weights[12][79] = 16'sd-37;
        fc1_weights[12][80] = 16'sd-52;
        fc1_weights[12][81] = 16'sd-2;
        fc1_weights[12][82] = 16'sd41;
        fc1_weights[12][83] = 16'sd-37;
        fc1_weights[12][84] = 16'sd35;
        fc1_weights[12][85] = 16'sd7;
        fc1_weights[12][86] = 16'sd-36;
        fc1_weights[12][87] = 16'sd-89;
        fc1_weights[12][88] = 16'sd-34;
        fc1_weights[12][89] = 16'sd-31;
        fc1_weights[12][90] = 16'sd-64;
        fc1_weights[12][91] = 16'sd-68;
        fc1_weights[12][92] = 16'sd-15;
        fc1_weights[12][93] = 16'sd5;
        fc1_weights[12][94] = 16'sd-27;
        fc1_weights[12][95] = 16'sd-36;
        fc1_weights[12][96] = 16'sd11;
        fc1_weights[12][97] = 16'sd-85;
        fc1_weights[12][98] = 16'sd12;
        fc1_weights[12][99] = 16'sd-60;
        fc1_weights[12][100] = 16'sd-107;
        fc1_weights[12][101] = 16'sd13;
        fc1_weights[12][102] = 16'sd-38;
        fc1_weights[12][103] = 16'sd5;
        fc1_weights[12][104] = 16'sd38;
        fc1_weights[12][105] = 16'sd118;
        fc1_weights[12][106] = 16'sd22;
        fc1_weights[12][107] = 16'sd-59;
        fc1_weights[12][108] = 16'sd3;
        fc1_weights[12][109] = 16'sd39;
        fc1_weights[12][110] = 16'sd-5;
        fc1_weights[12][111] = 16'sd25;
        fc1_weights[12][112] = 16'sd-104;
        fc1_weights[12][113] = 16'sd-100;
        fc1_weights[12][114] = 16'sd70;
        fc1_weights[12][115] = 16'sd93;
        fc1_weights[12][116] = 16'sd3;
        fc1_weights[12][117] = 16'sd-73;
        fc1_weights[12][118] = 16'sd-29;
        fc1_weights[12][119] = 16'sd-80;
        fc1_weights[12][120] = 16'sd-98;
        fc1_weights[12][121] = 16'sd21;
        fc1_weights[12][122] = 16'sd-39;
        fc1_weights[12][123] = 16'sd-80;
        fc1_weights[12][124] = 16'sd-13;
        fc1_weights[12][125] = 16'sd0;
        fc1_weights[12][126] = 16'sd5;
        fc1_weights[12][127] = 16'sd29;
        fc1_weights[12][128] = 16'sd14;
        fc1_weights[12][129] = 16'sd51;
        fc1_weights[12][130] = 16'sd0;
        fc1_weights[12][131] = 16'sd17;
        fc1_weights[12][132] = 16'sd3;
        fc1_weights[12][133] = 16'sd30;
        fc1_weights[12][134] = 16'sd37;
        fc1_weights[12][135] = 16'sd34;
        fc1_weights[12][136] = 16'sd5;
        fc1_weights[12][137] = 16'sd3;
        fc1_weights[12][138] = 16'sd56;
        fc1_weights[12][139] = 16'sd63;
        fc1_weights[12][140] = 16'sd52;
        fc1_weights[12][141] = 16'sd65;
        fc1_weights[12][142] = 16'sd-63;
        fc1_weights[12][143] = 16'sd53;
        fc1_weights[12][144] = 16'sd-5;
        fc1_weights[12][145] = 16'sd49;
        fc1_weights[12][146] = 16'sd29;
        fc1_weights[12][147] = 16'sd-62;
        fc1_weights[12][148] = 16'sd-65;
        fc1_weights[12][149] = 16'sd-60;
        fc1_weights[12][150] = 16'sd20;
        fc1_weights[12][151] = 16'sd-13;
        fc1_weights[12][152] = 16'sd12;
        fc1_weights[12][153] = 16'sd-34;
        fc1_weights[12][154] = 16'sd-37;
        fc1_weights[12][155] = 16'sd-42;
        fc1_weights[12][156] = 16'sd-126;
        fc1_weights[12][157] = 16'sd-133;
        fc1_weights[12][158] = 16'sd12;
        fc1_weights[12][159] = 16'sd-10;
        fc1_weights[12][160] = 16'sd16;
        fc1_weights[12][161] = 16'sd-4;
        fc1_weights[12][162] = 16'sd-21;
        fc1_weights[12][163] = 16'sd4;
        fc1_weights[12][164] = 16'sd32;
        fc1_weights[12][165] = 16'sd3;
        fc1_weights[12][166] = 16'sd37;
        fc1_weights[12][167] = 16'sd2;
        fc1_weights[12][168] = 16'sd62;
        fc1_weights[12][169] = 16'sd7;
        fc1_weights[12][170] = 16'sd-69;
        fc1_weights[12][171] = 16'sd61;
        fc1_weights[12][172] = 16'sd16;
        fc1_weights[12][173] = 16'sd1;
        fc1_weights[12][174] = 16'sd40;
        fc1_weights[12][175] = 16'sd5;
        fc1_weights[12][176] = 16'sd-28;
        fc1_weights[12][177] = 16'sd-104;
        fc1_weights[12][178] = 16'sd-20;
        fc1_weights[12][179] = 16'sd35;
        fc1_weights[12][180] = 16'sd-40;
        fc1_weights[12][181] = 16'sd68;
        fc1_weights[12][182] = 16'sd18;
        fc1_weights[12][183] = 16'sd43;
        fc1_weights[12][184] = 16'sd87;
        fc1_weights[12][185] = 16'sd-11;
        fc1_weights[12][186] = 16'sd37;
        fc1_weights[12][187] = 16'sd45;
        fc1_weights[12][188] = 16'sd51;
        fc1_weights[12][189] = 16'sd41;
        fc1_weights[12][190] = 16'sd3;
        fc1_weights[12][191] = 16'sd16;
        fc1_weights[12][192] = 16'sd40;
        fc1_weights[12][193] = 16'sd45;
        fc1_weights[12][194] = 16'sd-43;
        fc1_weights[12][195] = 16'sd-71;
        fc1_weights[12][196] = 16'sd1;
        fc1_weights[12][197] = 16'sd-27;
        fc1_weights[12][198] = 16'sd75;
        fc1_weights[12][199] = 16'sd-34;
        fc1_weights[12][200] = 16'sd15;
        fc1_weights[12][201] = 16'sd12;
        fc1_weights[12][202] = 16'sd-9;
        fc1_weights[12][203] = 16'sd-114;
        fc1_weights[12][204] = 16'sd-14;
        fc1_weights[12][205] = 16'sd16;
        fc1_weights[12][206] = 16'sd23;
        fc1_weights[12][207] = 16'sd57;
        fc1_weights[13][0] = 16'sd-26;
        fc1_weights[13][1] = 16'sd4;
        fc1_weights[13][2] = 16'sd19;
        fc1_weights[13][3] = 16'sd7;
        fc1_weights[13][4] = 16'sd2;
        fc1_weights[13][5] = 16'sd-11;
        fc1_weights[13][6] = 16'sd2;
        fc1_weights[13][7] = 16'sd18;
        fc1_weights[13][8] = 16'sd10;
        fc1_weights[13][9] = 16'sd23;
        fc1_weights[13][10] = 16'sd-9;
        fc1_weights[13][11] = 16'sd19;
        fc1_weights[13][12] = 16'sd7;
        fc1_weights[13][13] = 16'sd-22;
        fc1_weights[13][14] = 16'sd-27;
        fc1_weights[13][15] = 16'sd-18;
        fc1_weights[13][16] = 16'sd-7;
        fc1_weights[13][17] = 16'sd15;
        fc1_weights[13][18] = 16'sd6;
        fc1_weights[13][19] = 16'sd-5;
        fc1_weights[13][20] = 16'sd61;
        fc1_weights[13][21] = 16'sd22;
        fc1_weights[13][22] = 16'sd22;
        fc1_weights[13][23] = 16'sd19;
        fc1_weights[13][24] = 16'sd29;
        fc1_weights[13][25] = 16'sd7;
        fc1_weights[13][26] = 16'sd-36;
        fc1_weights[13][27] = 16'sd-18;
        fc1_weights[13][28] = 16'sd5;
        fc1_weights[13][29] = 16'sd-20;
        fc1_weights[13][30] = 16'sd-4;
        fc1_weights[13][31] = 16'sd5;
        fc1_weights[13][32] = 16'sd-16;
        fc1_weights[13][33] = 16'sd-7;
        fc1_weights[13][34] = 16'sd-28;
        fc1_weights[13][35] = 16'sd-13;
        fc1_weights[13][36] = 16'sd17;
        fc1_weights[13][37] = 16'sd9;
        fc1_weights[13][38] = 16'sd0;
        fc1_weights[13][39] = 16'sd10;
        fc1_weights[13][40] = 16'sd8;
        fc1_weights[13][41] = 16'sd-40;
        fc1_weights[13][42] = 16'sd27;
        fc1_weights[13][43] = 16'sd21;
        fc1_weights[13][44] = 16'sd-28;
        fc1_weights[13][45] = 16'sd-21;
        fc1_weights[13][46] = 16'sd-1;
        fc1_weights[13][47] = 16'sd19;
        fc1_weights[13][48] = 16'sd-9;
        fc1_weights[13][49] = 16'sd-4;
        fc1_weights[13][50] = 16'sd1;
        fc1_weights[13][51] = 16'sd-25;
        fc1_weights[13][52] = 16'sd-25;
        fc1_weights[13][53] = 16'sd-8;
        fc1_weights[13][54] = 16'sd3;
        fc1_weights[13][55] = 16'sd-1;
        fc1_weights[13][56] = 16'sd16;
        fc1_weights[13][57] = 16'sd22;
        fc1_weights[13][58] = 16'sd1;
        fc1_weights[13][59] = 16'sd10;
        fc1_weights[13][60] = 16'sd0;
        fc1_weights[13][61] = 16'sd21;
        fc1_weights[13][62] = 16'sd-17;
        fc1_weights[13][63] = 16'sd13;
        fc1_weights[13][64] = 16'sd-5;
        fc1_weights[13][65] = 16'sd-31;
        fc1_weights[13][66] = 16'sd-17;
        fc1_weights[13][67] = 16'sd6;
        fc1_weights[13][68] = 16'sd-18;
        fc1_weights[13][69] = 16'sd-10;
        fc1_weights[13][70] = 16'sd-23;
        fc1_weights[13][71] = 16'sd29;
        fc1_weights[13][72] = 16'sd31;
        fc1_weights[13][73] = 16'sd2;
        fc1_weights[13][74] = 16'sd16;
        fc1_weights[13][75] = 16'sd8;
        fc1_weights[13][76] = 16'sd-6;
        fc1_weights[13][77] = 16'sd15;
        fc1_weights[13][78] = 16'sd19;
        fc1_weights[13][79] = 16'sd14;
        fc1_weights[13][80] = 16'sd8;
        fc1_weights[13][81] = 16'sd-17;
        fc1_weights[13][82] = 16'sd-15;
        fc1_weights[13][83] = 16'sd12;
        fc1_weights[13][84] = 16'sd12;
        fc1_weights[13][85] = 16'sd7;
        fc1_weights[13][86] = 16'sd20;
        fc1_weights[13][87] = 16'sd13;
        fc1_weights[13][88] = 16'sd-42;
        fc1_weights[13][89] = 16'sd-3;
        fc1_weights[13][90] = 16'sd13;
        fc1_weights[13][91] = 16'sd-18;
        fc1_weights[13][92] = 16'sd12;
        fc1_weights[13][93] = 16'sd-14;
        fc1_weights[13][94] = 16'sd-18;
        fc1_weights[13][95] = 16'sd-11;
        fc1_weights[13][96] = 16'sd-30;
        fc1_weights[13][97] = 16'sd-28;
        fc1_weights[13][98] = 16'sd-15;
        fc1_weights[13][99] = 16'sd-13;
        fc1_weights[13][100] = 16'sd28;
        fc1_weights[13][101] = 16'sd28;
        fc1_weights[13][102] = 16'sd41;
        fc1_weights[13][103] = 16'sd3;
        fc1_weights[13][104] = 16'sd6;
        fc1_weights[13][105] = 16'sd-50;
        fc1_weights[13][106] = 16'sd2;
        fc1_weights[13][107] = 16'sd-15;
        fc1_weights[13][108] = 16'sd-28;
        fc1_weights[13][109] = 16'sd-7;
        fc1_weights[13][110] = 16'sd39;
        fc1_weights[13][111] = 16'sd20;
        fc1_weights[13][112] = 16'sd-7;
        fc1_weights[13][113] = 16'sd-12;
        fc1_weights[13][114] = 16'sd-21;
        fc1_weights[13][115] = 16'sd-1;
        fc1_weights[13][116] = 16'sd10;
        fc1_weights[13][117] = 16'sd-2;
        fc1_weights[13][118] = 16'sd25;
        fc1_weights[13][119] = 16'sd20;
        fc1_weights[13][120] = 16'sd-6;
        fc1_weights[13][121] = 16'sd-10;
        fc1_weights[13][122] = 16'sd-29;
        fc1_weights[13][123] = 16'sd-6;
        fc1_weights[13][124] = 16'sd12;
        fc1_weights[13][125] = 16'sd28;
        fc1_weights[13][126] = 16'sd-20;
        fc1_weights[13][127] = 16'sd9;
        fc1_weights[13][128] = 16'sd20;
        fc1_weights[13][129] = 16'sd-15;
        fc1_weights[13][130] = 16'sd32;
        fc1_weights[13][131] = 16'sd21;
        fc1_weights[13][132] = 16'sd14;
        fc1_weights[13][133] = 16'sd2;
        fc1_weights[13][134] = 16'sd-29;
        fc1_weights[13][135] = 16'sd-14;
        fc1_weights[13][136] = 16'sd27;
        fc1_weights[13][137] = 16'sd8;
        fc1_weights[13][138] = 16'sd-22;
        fc1_weights[13][139] = 16'sd-34;
        fc1_weights[13][140] = 16'sd-23;
        fc1_weights[13][141] = 16'sd-12;
        fc1_weights[13][142] = 16'sd-23;
        fc1_weights[13][143] = 16'sd-26;
        fc1_weights[13][144] = 16'sd-6;
        fc1_weights[13][145] = 16'sd9;
        fc1_weights[13][146] = 16'sd29;
        fc1_weights[13][147] = 16'sd28;
        fc1_weights[13][148] = 16'sd-5;
        fc1_weights[13][149] = 16'sd-23;
        fc1_weights[13][150] = 16'sd-10;
        fc1_weights[13][151] = 16'sd-2;
        fc1_weights[13][152] = 16'sd-10;
        fc1_weights[13][153] = 16'sd39;
        fc1_weights[13][154] = 16'sd-4;
        fc1_weights[13][155] = 16'sd20;
        fc1_weights[13][156] = 16'sd4;
        fc1_weights[13][157] = 16'sd-6;
        fc1_weights[13][158] = 16'sd8;
        fc1_weights[13][159] = 16'sd0;
        fc1_weights[13][160] = 16'sd-20;
        fc1_weights[13][161] = 16'sd14;
        fc1_weights[13][162] = 16'sd-4;
        fc1_weights[13][163] = 16'sd-13;
        fc1_weights[13][164] = 16'sd-2;
        fc1_weights[13][165] = 16'sd-24;
        fc1_weights[13][166] = 16'sd5;
        fc1_weights[13][167] = 16'sd-9;
        fc1_weights[13][168] = 16'sd-10;
        fc1_weights[13][169] = 16'sd9;
        fc1_weights[13][170] = 16'sd15;
        fc1_weights[13][171] = 16'sd18;
        fc1_weights[13][172] = 16'sd-9;
        fc1_weights[13][173] = 16'sd30;
        fc1_weights[13][174] = 16'sd31;
        fc1_weights[13][175] = 16'sd36;
        fc1_weights[13][176] = 16'sd22;
        fc1_weights[13][177] = 16'sd-14;
        fc1_weights[13][178] = 16'sd2;
        fc1_weights[13][179] = 16'sd10;
        fc1_weights[13][180] = 16'sd-19;
        fc1_weights[13][181] = 16'sd-22;
        fc1_weights[13][182] = 16'sd-11;
        fc1_weights[13][183] = 16'sd-12;
        fc1_weights[13][184] = 16'sd-20;
        fc1_weights[13][185] = 16'sd-7;
        fc1_weights[13][186] = 16'sd-48;
        fc1_weights[13][187] = 16'sd-11;
        fc1_weights[13][188] = 16'sd-7;
        fc1_weights[13][189] = 16'sd-15;
        fc1_weights[13][190] = 16'sd-14;
        fc1_weights[13][191] = 16'sd-13;
        fc1_weights[13][192] = 16'sd4;
        fc1_weights[13][193] = 16'sd2;
        fc1_weights[13][194] = 16'sd0;
        fc1_weights[13][195] = 16'sd-9;
        fc1_weights[13][196] = 16'sd14;
        fc1_weights[13][197] = 16'sd4;
        fc1_weights[13][198] = 16'sd10;
        fc1_weights[13][199] = 16'sd16;
        fc1_weights[13][200] = 16'sd23;
        fc1_weights[13][201] = 16'sd27;
        fc1_weights[13][202] = 16'sd40;
        fc1_weights[13][203] = 16'sd0;
        fc1_weights[13][204] = 16'sd25;
        fc1_weights[13][205] = 16'sd-4;
        fc1_weights[13][206] = 16'sd4;
        fc1_weights[13][207] = 16'sd1;
        fc1_weights[14][0] = 16'sd27;
        fc1_weights[14][1] = 16'sd32;
        fc1_weights[14][2] = 16'sd-18;
        fc1_weights[14][3] = 16'sd-35;
        fc1_weights[14][4] = 16'sd-73;
        fc1_weights[14][5] = 16'sd6;
        fc1_weights[14][6] = 16'sd26;
        fc1_weights[14][7] = 16'sd33;
        fc1_weights[14][8] = 16'sd-22;
        fc1_weights[14][9] = 16'sd-54;
        fc1_weights[14][10] = 16'sd-38;
        fc1_weights[14][11] = 16'sd-88;
        fc1_weights[14][12] = 16'sd-106;
        fc1_weights[14][13] = 16'sd-7;
        fc1_weights[14][14] = 16'sd90;
        fc1_weights[14][15] = 16'sd104;
        fc1_weights[14][16] = 16'sd119;
        fc1_weights[14][17] = 16'sd46;
        fc1_weights[14][18] = 16'sd27;
        fc1_weights[14][19] = 16'sd-26;
        fc1_weights[14][20] = 16'sd56;
        fc1_weights[14][21] = 16'sd15;
        fc1_weights[14][22] = 16'sd51;
        fc1_weights[14][23] = 16'sd35;
        fc1_weights[14][24] = 16'sd12;
        fc1_weights[14][25] = 16'sd22;
        fc1_weights[14][26] = 16'sd-6;
        fc1_weights[14][27] = 16'sd6;
        fc1_weights[14][28] = 16'sd-8;
        fc1_weights[14][29] = 16'sd-31;
        fc1_weights[14][30] = 16'sd-11;
        fc1_weights[14][31] = 16'sd26;
        fc1_weights[14][32] = 16'sd36;
        fc1_weights[14][33] = 16'sd-47;
        fc1_weights[14][34] = 16'sd-15;
        fc1_weights[14][35] = 16'sd-23;
        fc1_weights[14][36] = 16'sd-17;
        fc1_weights[14][37] = 16'sd-59;
        fc1_weights[14][38] = 16'sd-7;
        fc1_weights[14][39] = 16'sd5;
        fc1_weights[14][40] = 16'sd115;
        fc1_weights[14][41] = 16'sd120;
        fc1_weights[14][42] = 16'sd31;
        fc1_weights[14][43] = 16'sd27;
        fc1_weights[14][44] = 16'sd24;
        fc1_weights[14][45] = 16'sd-62;
        fc1_weights[14][46] = 16'sd-33;
        fc1_weights[14][47] = 16'sd-64;
        fc1_weights[14][48] = 16'sd-35;
        fc1_weights[14][49] = 16'sd-9;
        fc1_weights[14][50] = 16'sd5;
        fc1_weights[14][51] = 16'sd-59;
        fc1_weights[14][52] = 16'sd-28;
        fc1_weights[14][53] = 16'sd27;
        fc1_weights[14][54] = 16'sd-32;
        fc1_weights[14][55] = 16'sd-41;
        fc1_weights[14][56] = 16'sd11;
        fc1_weights[14][57] = 16'sd13;
        fc1_weights[14][58] = 16'sd50;
        fc1_weights[14][59] = 16'sd-10;
        fc1_weights[14][60] = 16'sd-37;
        fc1_weights[14][61] = 16'sd-6;
        fc1_weights[14][62] = 16'sd-35;
        fc1_weights[14][63] = 16'sd17;
        fc1_weights[14][64] = 16'sd38;
        fc1_weights[14][65] = 16'sd-47;
        fc1_weights[14][66] = 16'sd29;
        fc1_weights[14][67] = 16'sd74;
        fc1_weights[14][68] = 16'sd-19;
        fc1_weights[14][69] = 16'sd-1;
        fc1_weights[14][70] = 16'sd47;
        fc1_weights[14][71] = 16'sd6;
        fc1_weights[14][72] = 16'sd21;
        fc1_weights[14][73] = 16'sd-48;
        fc1_weights[14][74] = 16'sd-61;
        fc1_weights[14][75] = 16'sd-34;
        fc1_weights[14][76] = 16'sd-1;
        fc1_weights[14][77] = 16'sd-26;
        fc1_weights[14][78] = 16'sd-62;
        fc1_weights[14][79] = 16'sd24;
        fc1_weights[14][80] = 16'sd4;
        fc1_weights[14][81] = 16'sd-24;
        fc1_weights[14][82] = 16'sd-64;
        fc1_weights[14][83] = 16'sd-30;
        fc1_weights[14][84] = 16'sd34;
        fc1_weights[14][85] = 16'sd-25;
        fc1_weights[14][86] = 16'sd-18;
        fc1_weights[14][87] = 16'sd4;
        fc1_weights[14][88] = 16'sd-39;
        fc1_weights[14][89] = 16'sd46;
        fc1_weights[14][90] = 16'sd73;
        fc1_weights[14][91] = 16'sd82;
        fc1_weights[14][92] = 16'sd39;
        fc1_weights[14][93] = 16'sd122;
        fc1_weights[14][94] = 16'sd53;
        fc1_weights[14][95] = 16'sd20;
        fc1_weights[14][96] = 16'sd14;
        fc1_weights[14][97] = 16'sd14;
        fc1_weights[14][98] = 16'sd20;
        fc1_weights[14][99] = 16'sd-3;
        fc1_weights[14][100] = 16'sd-33;
        fc1_weights[14][101] = 16'sd-6;
        fc1_weights[14][102] = 16'sd-24;
        fc1_weights[14][103] = 16'sd-43;
        fc1_weights[14][104] = 16'sd-37;
        fc1_weights[14][105] = 16'sd-41;
        fc1_weights[14][106] = 16'sd-22;
        fc1_weights[14][107] = 16'sd-74;
        fc1_weights[14][108] = 16'sd32;
        fc1_weights[14][109] = 16'sd29;
        fc1_weights[14][110] = 16'sd37;
        fc1_weights[14][111] = 16'sd-37;
        fc1_weights[14][112] = 16'sd-20;
        fc1_weights[14][113] = 16'sd-28;
        fc1_weights[14][114] = 16'sd12;
        fc1_weights[14][115] = 16'sd-25;
        fc1_weights[14][116] = 16'sd-15;
        fc1_weights[14][117] = 16'sd-16;
        fc1_weights[14][118] = 16'sd-14;
        fc1_weights[14][119] = 16'sd27;
        fc1_weights[14][120] = 16'sd-1;
        fc1_weights[14][121] = 16'sd6;
        fc1_weights[14][122] = 16'sd-17;
        fc1_weights[14][123] = 16'sd-81;
        fc1_weights[14][124] = 16'sd-65;
        fc1_weights[14][125] = 16'sd-56;
        fc1_weights[14][126] = 16'sd-78;
        fc1_weights[14][127] = 16'sd-36;
        fc1_weights[14][128] = 16'sd-45;
        fc1_weights[14][129] = 16'sd-109;
        fc1_weights[14][130] = 16'sd-18;
        fc1_weights[14][131] = 16'sd-15;
        fc1_weights[14][132] = 16'sd-29;
        fc1_weights[14][133] = 16'sd3;
        fc1_weights[14][134] = 16'sd53;
        fc1_weights[14][135] = 16'sd40;
        fc1_weights[14][136] = 16'sd14;
        fc1_weights[14][137] = 16'sd-25;
        fc1_weights[14][138] = 16'sd-16;
        fc1_weights[14][139] = 16'sd24;
        fc1_weights[14][140] = 16'sd12;
        fc1_weights[14][141] = 16'sd38;
        fc1_weights[14][142] = 16'sd49;
        fc1_weights[14][143] = 16'sd30;
        fc1_weights[14][144] = 16'sd11;
        fc1_weights[14][145] = 16'sd-8;
        fc1_weights[14][146] = 16'sd9;
        fc1_weights[14][147] = 16'sd63;
        fc1_weights[14][148] = 16'sd-15;
        fc1_weights[14][149] = 16'sd-41;
        fc1_weights[14][150] = 16'sd-14;
        fc1_weights[14][151] = 16'sd-34;
        fc1_weights[14][152] = 16'sd30;
        fc1_weights[14][153] = 16'sd-8;
        fc1_weights[14][154] = 16'sd10;
        fc1_weights[14][155] = 16'sd7;
        fc1_weights[14][156] = 16'sd12;
        fc1_weights[14][157] = 16'sd-6;
        fc1_weights[14][158] = 16'sd-13;
        fc1_weights[14][159] = 16'sd-99;
        fc1_weights[14][160] = 16'sd-37;
        fc1_weights[14][161] = 16'sd-23;
        fc1_weights[14][162] = 16'sd-37;
        fc1_weights[14][163] = 16'sd-15;
        fc1_weights[14][164] = 16'sd-62;
        fc1_weights[14][165] = 16'sd23;
        fc1_weights[14][166] = 16'sd10;
        fc1_weights[14][167] = 16'sd33;
        fc1_weights[14][168] = 16'sd-10;
        fc1_weights[14][169] = 16'sd26;
        fc1_weights[14][170] = 16'sd47;
        fc1_weights[14][171] = 16'sd-3;
        fc1_weights[14][172] = 16'sd17;
        fc1_weights[14][173] = 16'sd22;
        fc1_weights[14][174] = 16'sd37;
        fc1_weights[14][175] = 16'sd17;
        fc1_weights[14][176] = 16'sd11;
        fc1_weights[14][177] = 16'sd-32;
        fc1_weights[14][178] = 16'sd-31;
        fc1_weights[14][179] = 16'sd15;
        fc1_weights[14][180] = 16'sd-18;
        fc1_weights[14][181] = 16'sd27;
        fc1_weights[14][182] = 16'sd1;
        fc1_weights[14][183] = 16'sd3;
        fc1_weights[14][184] = 16'sd-15;
        fc1_weights[14][185] = 16'sd-52;
        fc1_weights[14][186] = 16'sd-54;
        fc1_weights[14][187] = 16'sd-62;
        fc1_weights[14][188] = 16'sd-103;
        fc1_weights[14][189] = 16'sd-80;
        fc1_weights[14][190] = 16'sd15;
        fc1_weights[14][191] = 16'sd11;
        fc1_weights[14][192] = 16'sd-23;
        fc1_weights[14][193] = 16'sd-12;
        fc1_weights[14][194] = 16'sd12;
        fc1_weights[14][195] = 16'sd35;
        fc1_weights[14][196] = 16'sd30;
        fc1_weights[14][197] = 16'sd-3;
        fc1_weights[14][198] = 16'sd-15;
        fc1_weights[14][199] = 16'sd39;
        fc1_weights[14][200] = 16'sd19;
        fc1_weights[14][201] = 16'sd-26;
        fc1_weights[14][202] = 16'sd-26;
        fc1_weights[14][203] = 16'sd44;
        fc1_weights[14][204] = 16'sd0;
        fc1_weights[14][205] = 16'sd21;
        fc1_weights[14][206] = 16'sd22;
        fc1_weights[14][207] = 16'sd39;
        fc1_weights[15][0] = 16'sd-5;
        fc1_weights[15][1] = 16'sd-1;
        fc1_weights[15][2] = 16'sd-14;
        fc1_weights[15][3] = 16'sd5;
        fc1_weights[15][4] = 16'sd-33;
        fc1_weights[15][5] = 16'sd-34;
        fc1_weights[15][6] = 16'sd-65;
        fc1_weights[15][7] = 16'sd-38;
        fc1_weights[15][8] = 16'sd-41;
        fc1_weights[15][9] = 16'sd-22;
        fc1_weights[15][10] = 16'sd15;
        fc1_weights[15][11] = 16'sd-14;
        fc1_weights[15][12] = 16'sd-3;
        fc1_weights[15][13] = 16'sd-67;
        fc1_weights[15][14] = 16'sd-71;
        fc1_weights[15][15] = 16'sd-3;
        fc1_weights[15][16] = 16'sd-15;
        fc1_weights[15][17] = 16'sd-15;
        fc1_weights[15][18] = 16'sd28;
        fc1_weights[15][19] = 16'sd42;
        fc1_weights[15][20] = 16'sd33;
        fc1_weights[15][21] = 16'sd55;
        fc1_weights[15][22] = 16'sd30;
        fc1_weights[15][23] = 16'sd6;
        fc1_weights[15][24] = 16'sd23;
        fc1_weights[15][25] = 16'sd11;
        fc1_weights[15][26] = 16'sd-4;
        fc1_weights[15][27] = 16'sd-5;
        fc1_weights[15][28] = 16'sd8;
        fc1_weights[15][29] = 16'sd-7;
        fc1_weights[15][30] = 16'sd-46;
        fc1_weights[15][31] = 16'sd-18;
        fc1_weights[15][32] = 16'sd-45;
        fc1_weights[15][33] = 16'sd-19;
        fc1_weights[15][34] = 16'sd-48;
        fc1_weights[15][35] = 16'sd-23;
        fc1_weights[15][36] = 16'sd43;
        fc1_weights[15][37] = 16'sd-13;
        fc1_weights[15][38] = 16'sd-6;
        fc1_weights[15][39] = 16'sd-47;
        fc1_weights[15][40] = 16'sd-5;
        fc1_weights[15][41] = 16'sd-35;
        fc1_weights[15][42] = 16'sd7;
        fc1_weights[15][43] = 16'sd87;
        fc1_weights[15][44] = 16'sd30;
        fc1_weights[15][45] = 16'sd15;
        fc1_weights[15][46] = 16'sd2;
        fc1_weights[15][47] = 16'sd51;
        fc1_weights[15][48] = 16'sd54;
        fc1_weights[15][49] = 16'sd13;
        fc1_weights[15][50] = 16'sd3;
        fc1_weights[15][51] = 16'sd-19;
        fc1_weights[15][52] = 16'sd28;
        fc1_weights[15][53] = 16'sd42;
        fc1_weights[15][54] = 16'sd13;
        fc1_weights[15][55] = 16'sd9;
        fc1_weights[15][56] = 16'sd-16;
        fc1_weights[15][57] = 16'sd-15;
        fc1_weights[15][58] = 16'sd-43;
        fc1_weights[15][59] = 16'sd-35;
        fc1_weights[15][60] = 16'sd-16;
        fc1_weights[15][61] = 16'sd-12;
        fc1_weights[15][62] = 16'sd0;
        fc1_weights[15][63] = 16'sd8;
        fc1_weights[15][64] = 16'sd2;
        fc1_weights[15][65] = 16'sd-43;
        fc1_weights[15][66] = 16'sd25;
        fc1_weights[15][67] = 16'sd23;
        fc1_weights[15][68] = 16'sd37;
        fc1_weights[15][69] = 16'sd44;
        fc1_weights[15][70] = 16'sd14;
        fc1_weights[15][71] = 16'sd-7;
        fc1_weights[15][72] = 16'sd-4;
        fc1_weights[15][73] = 16'sd-39;
        fc1_weights[15][74] = 16'sd-21;
        fc1_weights[15][75] = 16'sd29;
        fc1_weights[15][76] = 16'sd-1;
        fc1_weights[15][77] = 16'sd-1;
        fc1_weights[15][78] = 16'sd50;
        fc1_weights[15][79] = 16'sd34;
        fc1_weights[15][80] = 16'sd-2;
        fc1_weights[15][81] = 16'sd-30;
        fc1_weights[15][82] = 16'sd12;
        fc1_weights[15][83] = 16'sd-18;
        fc1_weights[15][84] = 16'sd17;
        fc1_weights[15][85] = 16'sd1;
        fc1_weights[15][86] = 16'sd7;
        fc1_weights[15][87] = 16'sd-17;
        fc1_weights[15][88] = 16'sd-14;
        fc1_weights[15][89] = 16'sd38;
        fc1_weights[15][90] = 16'sd19;
        fc1_weights[15][91] = 16'sd49;
        fc1_weights[15][92] = 16'sd82;
        fc1_weights[15][93] = 16'sd66;
        fc1_weights[15][94] = 16'sd19;
        fc1_weights[15][95] = 16'sd-1;
        fc1_weights[15][96] = 16'sd-36;
        fc1_weights[15][97] = 16'sd-29;
        fc1_weights[15][98] = 16'sd-12;
        fc1_weights[15][99] = 16'sd-14;
        fc1_weights[15][100] = 16'sd-31;
        fc1_weights[15][101] = 16'sd-1;
        fc1_weights[15][102] = 16'sd19;
        fc1_weights[15][103] = 16'sd13;
        fc1_weights[15][104] = 16'sd25;
        fc1_weights[15][105] = 16'sd5;
        fc1_weights[15][106] = 16'sd32;
        fc1_weights[15][107] = 16'sd17;
        fc1_weights[15][108] = 16'sd12;
        fc1_weights[15][109] = 16'sd-21;
        fc1_weights[15][110] = 16'sd35;
        fc1_weights[15][111] = 16'sd1;
        fc1_weights[15][112] = 16'sd12;
        fc1_weights[15][113] = 16'sd22;
        fc1_weights[15][114] = 16'sd2;
        fc1_weights[15][115] = 16'sd7;
        fc1_weights[15][116] = 16'sd3;
        fc1_weights[15][117] = 16'sd22;
        fc1_weights[15][118] = 16'sd-3;
        fc1_weights[15][119] = 16'sd23;
        fc1_weights[15][120] = 16'sd-27;
        fc1_weights[15][121] = 16'sd20;
        fc1_weights[15][122] = 16'sd-14;
        fc1_weights[15][123] = 16'sd1;
        fc1_weights[15][124] = 16'sd5;
        fc1_weights[15][125] = 16'sd3;
        fc1_weights[15][126] = 16'sd-54;
        fc1_weights[15][127] = 16'sd-36;
        fc1_weights[15][128] = 16'sd-23;
        fc1_weights[15][129] = 16'sd-41;
        fc1_weights[15][130] = 16'sd7;
        fc1_weights[15][131] = 16'sd-32;
        fc1_weights[15][132] = 16'sd-1;
        fc1_weights[15][133] = 16'sd-27;
        fc1_weights[15][134] = 16'sd-23;
        fc1_weights[15][135] = 16'sd11;
        fc1_weights[15][136] = 16'sd5;
        fc1_weights[15][137] = 16'sd41;
        fc1_weights[15][138] = 16'sd15;
        fc1_weights[15][139] = 16'sd19;
        fc1_weights[15][140] = 16'sd-11;
        fc1_weights[15][141] = 16'sd2;
        fc1_weights[15][142] = 16'sd-8;
        fc1_weights[15][143] = 16'sd-26;
        fc1_weights[15][144] = 16'sd-19;
        fc1_weights[15][145] = 16'sd-4;
        fc1_weights[15][146] = 16'sd72;
        fc1_weights[15][147] = 16'sd41;
        fc1_weights[15][148] = 16'sd37;
        fc1_weights[15][149] = 16'sd8;
        fc1_weights[15][150] = 16'sd1;
        fc1_weights[15][151] = 16'sd-16;
        fc1_weights[15][152] = 16'sd-8;
        fc1_weights[15][153] = 16'sd8;
        fc1_weights[15][154] = 16'sd0;
        fc1_weights[15][155] = 16'sd-41;
        fc1_weights[15][156] = 16'sd37;
        fc1_weights[15][157] = 16'sd18;
        fc1_weights[15][158] = 16'sd7;
        fc1_weights[15][159] = 16'sd13;
        fc1_weights[15][160] = 16'sd-10;
        fc1_weights[15][161] = 16'sd11;
        fc1_weights[15][162] = 16'sd27;
        fc1_weights[15][163] = 16'sd8;
        fc1_weights[15][164] = 16'sd32;
        fc1_weights[15][165] = 16'sd-16;
        fc1_weights[15][166] = 16'sd-5;
        fc1_weights[15][167] = 16'sd2;
        fc1_weights[15][168] = 16'sd14;
        fc1_weights[15][169] = 16'sd-6;
        fc1_weights[15][170] = 16'sd-4;
        fc1_weights[15][171] = 16'sd23;
        fc1_weights[15][172] = 16'sd15;
        fc1_weights[15][173] = 16'sd43;
        fc1_weights[15][174] = 16'sd35;
        fc1_weights[15][175] = 16'sd28;
        fc1_weights[15][176] = 16'sd-35;
        fc1_weights[15][177] = 16'sd33;
        fc1_weights[15][178] = 16'sd13;
        fc1_weights[15][179] = 16'sd-22;
        fc1_weights[15][180] = 16'sd-8;
        fc1_weights[15][181] = 16'sd9;
        fc1_weights[15][182] = 16'sd17;
        fc1_weights[15][183] = 16'sd2;
        fc1_weights[15][184] = 16'sd-15;
        fc1_weights[15][185] = 16'sd25;
        fc1_weights[15][186] = 16'sd40;
        fc1_weights[15][187] = 16'sd28;
        fc1_weights[15][188] = 16'sd7;
        fc1_weights[15][189] = 16'sd8;
        fc1_weights[15][190] = 16'sd12;
        fc1_weights[15][191] = 16'sd14;
        fc1_weights[15][192] = 16'sd-31;
        fc1_weights[15][193] = 16'sd-16;
        fc1_weights[15][194] = 16'sd-4;
        fc1_weights[15][195] = 16'sd-13;
        fc1_weights[15][196] = 16'sd-10;
        fc1_weights[15][197] = 16'sd25;
        fc1_weights[15][198] = 16'sd21;
        fc1_weights[15][199] = 16'sd36;
        fc1_weights[15][200] = 16'sd37;
        fc1_weights[15][201] = 16'sd71;
        fc1_weights[15][202] = 16'sd6;
        fc1_weights[15][203] = 16'sd32;
        fc1_weights[15][204] = 16'sd24;
        fc1_weights[15][205] = 16'sd46;
        fc1_weights[15][206] = 16'sd-3;
        fc1_weights[15][207] = 16'sd-16;
        fc1_weights[16][0] = 16'sd-12;
        fc1_weights[16][1] = 16'sd8;
        fc1_weights[16][2] = 16'sd41;
        fc1_weights[16][3] = 16'sd34;
        fc1_weights[16][4] = 16'sd-16;
        fc1_weights[16][5] = 16'sd23;
        fc1_weights[16][6] = 16'sd4;
        fc1_weights[16][7] = 16'sd-37;
        fc1_weights[16][8] = 16'sd-4;
        fc1_weights[16][9] = 16'sd-52;
        fc1_weights[16][10] = 16'sd-48;
        fc1_weights[16][11] = 16'sd-29;
        fc1_weights[16][12] = 16'sd23;
        fc1_weights[16][13] = 16'sd8;
        fc1_weights[16][14] = 16'sd-17;
        fc1_weights[16][15] = 16'sd27;
        fc1_weights[16][16] = 16'sd16;
        fc1_weights[16][17] = 16'sd-16;
        fc1_weights[16][18] = 16'sd34;
        fc1_weights[16][19] = 16'sd-24;
        fc1_weights[16][20] = 16'sd-9;
        fc1_weights[16][21] = 16'sd12;
        fc1_weights[16][22] = 16'sd-13;
        fc1_weights[16][23] = 16'sd14;
        fc1_weights[16][24] = 16'sd18;
        fc1_weights[16][25] = 16'sd35;
        fc1_weights[16][26] = 16'sd-41;
        fc1_weights[16][27] = 16'sd-68;
        fc1_weights[16][28] = 16'sd-20;
        fc1_weights[16][29] = 16'sd31;
        fc1_weights[16][30] = 16'sd38;
        fc1_weights[16][31] = 16'sd-4;
        fc1_weights[16][32] = 16'sd16;
        fc1_weights[16][33] = 16'sd-82;
        fc1_weights[16][34] = 16'sd2;
        fc1_weights[16][35] = 16'sd-12;
        fc1_weights[16][36] = 16'sd-3;
        fc1_weights[16][37] = 16'sd-68;
        fc1_weights[16][38] = 16'sd27;
        fc1_weights[16][39] = 16'sd17;
        fc1_weights[16][40] = 16'sd34;
        fc1_weights[16][41] = 16'sd58;
        fc1_weights[16][42] = 16'sd9;
        fc1_weights[16][43] = 16'sd-48;
        fc1_weights[16][44] = 16'sd-19;
        fc1_weights[16][45] = 16'sd-29;
        fc1_weights[16][46] = 16'sd-32;
        fc1_weights[16][47] = 16'sd1;
        fc1_weights[16][48] = 16'sd-50;
        fc1_weights[16][49] = 16'sd-19;
        fc1_weights[16][50] = 16'sd-50;
        fc1_weights[16][51] = 16'sd-42;
        fc1_weights[16][52] = 16'sd29;
        fc1_weights[16][53] = 16'sd13;
        fc1_weights[16][54] = 16'sd14;
        fc1_weights[16][55] = 16'sd-18;
        fc1_weights[16][56] = 16'sd65;
        fc1_weights[16][57] = 16'sd4;
        fc1_weights[16][58] = 16'sd33;
        fc1_weights[16][59] = 16'sd36;
        fc1_weights[16][60] = 16'sd74;
        fc1_weights[16][61] = 16'sd-7;
        fc1_weights[16][62] = 16'sd-35;
        fc1_weights[16][63] = 16'sd-15;
        fc1_weights[16][64] = 16'sd68;
        fc1_weights[16][65] = 16'sd31;
        fc1_weights[16][66] = 16'sd81;
        fc1_weights[16][67] = 16'sd34;
        fc1_weights[16][68] = 16'sd14;
        fc1_weights[16][69] = 16'sd-17;
        fc1_weights[16][70] = 16'sd20;
        fc1_weights[16][71] = 16'sd36;
        fc1_weights[16][72] = 16'sd-11;
        fc1_weights[16][73] = 16'sd18;
        fc1_weights[16][74] = 16'sd45;
        fc1_weights[16][75] = 16'sd-24;
        fc1_weights[16][76] = 16'sd-32;
        fc1_weights[16][77] = 16'sd14;
        fc1_weights[16][78] = 16'sd18;
        fc1_weights[16][79] = 16'sd10;
        fc1_weights[16][80] = 16'sd-5;
        fc1_weights[16][81] = 16'sd6;
        fc1_weights[16][82] = 16'sd19;
        fc1_weights[16][83] = 16'sd-10;
        fc1_weights[16][84] = 16'sd-10;
        fc1_weights[16][85] = 16'sd12;
        fc1_weights[16][86] = 16'sd48;
        fc1_weights[16][87] = 16'sd36;
        fc1_weights[16][88] = 16'sd-2;
        fc1_weights[16][89] = 16'sd0;
        fc1_weights[16][90] = 16'sd18;
        fc1_weights[16][91] = 16'sd74;
        fc1_weights[16][92] = 16'sd73;
        fc1_weights[16][93] = 16'sd11;
        fc1_weights[16][94] = 16'sd-13;
        fc1_weights[16][95] = 16'sd32;
        fc1_weights[16][96] = 16'sd34;
        fc1_weights[16][97] = 16'sd48;
        fc1_weights[16][98] = 16'sd35;
        fc1_weights[16][99] = 16'sd16;
        fc1_weights[16][100] = 16'sd24;
        fc1_weights[16][101] = 16'sd12;
        fc1_weights[16][102] = 16'sd-22;
        fc1_weights[16][103] = 16'sd11;
        fc1_weights[16][104] = 16'sd35;
        fc1_weights[16][105] = 16'sd6;
        fc1_weights[16][106] = 16'sd52;
        fc1_weights[16][107] = 16'sd13;
        fc1_weights[16][108] = 16'sd5;
        fc1_weights[16][109] = 16'sd15;
        fc1_weights[16][110] = 16'sd9;
        fc1_weights[16][111] = 16'sd1;
        fc1_weights[16][112] = 16'sd30;
        fc1_weights[16][113] = 16'sd-16;
        fc1_weights[16][114] = 16'sd-32;
        fc1_weights[16][115] = 16'sd-58;
        fc1_weights[16][116] = 16'sd29;
        fc1_weights[16][117] = 16'sd19;
        fc1_weights[16][118] = 16'sd17;
        fc1_weights[16][119] = 16'sd39;
        fc1_weights[16][120] = 16'sd15;
        fc1_weights[16][121] = 16'sd23;
        fc1_weights[16][122] = 16'sd31;
        fc1_weights[16][123] = 16'sd112;
        fc1_weights[16][124] = 16'sd5;
        fc1_weights[16][125] = 16'sd42;
        fc1_weights[16][126] = 16'sd20;
        fc1_weights[16][127] = 16'sd20;
        fc1_weights[16][128] = 16'sd23;
        fc1_weights[16][129] = 16'sd15;
        fc1_weights[16][130] = 16'sd-53;
        fc1_weights[16][131] = 16'sd-3;
        fc1_weights[16][132] = 16'sd-3;
        fc1_weights[16][133] = 16'sd14;
        fc1_weights[16][134] = 16'sd32;
        fc1_weights[16][135] = 16'sd45;
        fc1_weights[16][136] = 16'sd-32;
        fc1_weights[16][137] = 16'sd-30;
        fc1_weights[16][138] = 16'sd21;
        fc1_weights[16][139] = 16'sd-20;
        fc1_weights[16][140] = 16'sd-46;
        fc1_weights[16][141] = 16'sd-43;
        fc1_weights[16][142] = 16'sd25;
        fc1_weights[16][143] = 16'sd-21;
        fc1_weights[16][144] = 16'sd18;
        fc1_weights[16][145] = 16'sd-41;
        fc1_weights[16][146] = 16'sd-32;
        fc1_weights[16][147] = 16'sd-9;
        fc1_weights[16][148] = 16'sd-24;
        fc1_weights[16][149] = 16'sd-6;
        fc1_weights[16][150] = 16'sd22;
        fc1_weights[16][151] = 16'sd71;
        fc1_weights[16][152] = 16'sd-48;
        fc1_weights[16][153] = 16'sd-4;
        fc1_weights[16][154] = 16'sd4;
        fc1_weights[16][155] = 16'sd65;
        fc1_weights[16][156] = 16'sd1;
        fc1_weights[16][157] = 16'sd11;
        fc1_weights[16][158] = 16'sd-20;
        fc1_weights[16][159] = 16'sd-26;
        fc1_weights[16][160] = 16'sd-14;
        fc1_weights[16][161] = 16'sd15;
        fc1_weights[16][162] = 16'sd47;
        fc1_weights[16][163] = 16'sd-2;
        fc1_weights[16][164] = 16'sd-48;
        fc1_weights[16][165] = 16'sd-20;
        fc1_weights[16][166] = 16'sd-37;
        fc1_weights[16][167] = 16'sd0;
        fc1_weights[16][168] = 16'sd8;
        fc1_weights[16][169] = 16'sd10;
        fc1_weights[16][170] = 16'sd24;
        fc1_weights[16][171] = 16'sd-61;
        fc1_weights[16][172] = 16'sd-44;
        fc1_weights[16][173] = 16'sd-35;
        fc1_weights[16][174] = 16'sd-27;
        fc1_weights[16][175] = 16'sd-15;
        fc1_weights[16][176] = 16'sd-8;
        fc1_weights[16][177] = 16'sd19;
        fc1_weights[16][178] = 16'sd0;
        fc1_weights[16][179] = 16'sd59;
        fc1_weights[16][180] = 16'sd56;
        fc1_weights[16][181] = 16'sd55;
        fc1_weights[16][182] = 16'sd-14;
        fc1_weights[16][183] = 16'sd0;
        fc1_weights[16][184] = 16'sd10;
        fc1_weights[16][185] = 16'sd-5;
        fc1_weights[16][186] = 16'sd-25;
        fc1_weights[16][187] = 16'sd-30;
        fc1_weights[16][188] = 16'sd-18;
        fc1_weights[16][189] = 16'sd13;
        fc1_weights[16][190] = 16'sd37;
        fc1_weights[16][191] = 16'sd34;
        fc1_weights[16][192] = 16'sd47;
        fc1_weights[16][193] = 16'sd51;
        fc1_weights[16][194] = 16'sd34;
        fc1_weights[16][195] = 16'sd36;
        fc1_weights[16][196] = 16'sd14;
        fc1_weights[16][197] = 16'sd43;
        fc1_weights[16][198] = 16'sd-31;
        fc1_weights[16][199] = 16'sd-43;
        fc1_weights[16][200] = 16'sd-25;
        fc1_weights[16][201] = 16'sd-40;
        fc1_weights[16][202] = 16'sd-64;
        fc1_weights[16][203] = 16'sd16;
        fc1_weights[16][204] = 16'sd2;
        fc1_weights[16][205] = 16'sd-21;
        fc1_weights[16][206] = 16'sd-20;
        fc1_weights[16][207] = 16'sd45;
        fc1_weights[17][0] = 16'sd-10;
        fc1_weights[17][1] = 16'sd10;
        fc1_weights[17][2] = 16'sd21;
        fc1_weights[17][3] = 16'sd60;
        fc1_weights[17][4] = 16'sd-4;
        fc1_weights[17][5] = 16'sd-19;
        fc1_weights[17][6] = 16'sd4;
        fc1_weights[17][7] = 16'sd-14;
        fc1_weights[17][8] = 16'sd38;
        fc1_weights[17][9] = 16'sd43;
        fc1_weights[17][10] = 16'sd0;
        fc1_weights[17][11] = 16'sd55;
        fc1_weights[17][12] = 16'sd0;
        fc1_weights[17][13] = 16'sd54;
        fc1_weights[17][14] = 16'sd-34;
        fc1_weights[17][15] = 16'sd-86;
        fc1_weights[17][16] = 16'sd-72;
        fc1_weights[17][17] = 16'sd-36;
        fc1_weights[17][18] = 16'sd-77;
        fc1_weights[17][19] = 16'sd-33;
        fc1_weights[17][20] = 16'sd12;
        fc1_weights[17][21] = 16'sd-51;
        fc1_weights[17][22] = 16'sd18;
        fc1_weights[17][23] = 16'sd41;
        fc1_weights[17][24] = 16'sd35;
        fc1_weights[17][25] = 16'sd2;
        fc1_weights[17][26] = 16'sd-31;
        fc1_weights[17][27] = 16'sd-25;
        fc1_weights[17][28] = 16'sd43;
        fc1_weights[17][29] = 16'sd-13;
        fc1_weights[17][30] = 16'sd-6;
        fc1_weights[17][31] = 16'sd6;
        fc1_weights[17][32] = 16'sd2;
        fc1_weights[17][33] = 16'sd-35;
        fc1_weights[17][34] = 16'sd-66;
        fc1_weights[17][35] = 16'sd-8;
        fc1_weights[17][36] = 16'sd-13;
        fc1_weights[17][37] = 16'sd-16;
        fc1_weights[17][38] = 16'sd-13;
        fc1_weights[17][39] = 16'sd-16;
        fc1_weights[17][40] = 16'sd-9;
        fc1_weights[17][41] = 16'sd-70;
        fc1_weights[17][42] = 16'sd5;
        fc1_weights[17][43] = 16'sd-18;
        fc1_weights[17][44] = 16'sd-52;
        fc1_weights[17][45] = 16'sd-31;
        fc1_weights[17][46] = 16'sd-17;
        fc1_weights[17][47] = 16'sd21;
        fc1_weights[17][48] = 16'sd-31;
        fc1_weights[17][49] = 16'sd-17;
        fc1_weights[17][50] = 16'sd-27;
        fc1_weights[17][51] = 16'sd-38;
        fc1_weights[17][52] = 16'sd-37;
        fc1_weights[17][53] = 16'sd8;
        fc1_weights[17][54] = 16'sd9;
        fc1_weights[17][55] = 16'sd-71;
        fc1_weights[17][56] = 16'sd4;
        fc1_weights[17][57] = 16'sd5;
        fc1_weights[17][58] = 16'sd-19;
        fc1_weights[17][59] = 16'sd-33;
        fc1_weights[17][60] = 16'sd-51;
        fc1_weights[17][61] = 16'sd13;
        fc1_weights[17][62] = 16'sd-98;
        fc1_weights[17][63] = 16'sd-67;
        fc1_weights[17][64] = 16'sd-86;
        fc1_weights[17][65] = 16'sd-39;
        fc1_weights[17][66] = 16'sd-24;
        fc1_weights[17][67] = 16'sd-53;
        fc1_weights[17][68] = 16'sd-4;
        fc1_weights[17][69] = 16'sd-25;
        fc1_weights[17][70] = 16'sd-73;
        fc1_weights[17][71] = 16'sd-3;
        fc1_weights[17][72] = 16'sd37;
        fc1_weights[17][73] = 16'sd17;
        fc1_weights[17][74] = 16'sd12;
        fc1_weights[17][75] = 16'sd68;
        fc1_weights[17][76] = 16'sd20;
        fc1_weights[17][77] = 16'sd-15;
        fc1_weights[17][78] = 16'sd-43;
        fc1_weights[17][79] = 16'sd-4;
        fc1_weights[17][80] = 16'sd17;
        fc1_weights[17][81] = 16'sd24;
        fc1_weights[17][82] = 16'sd1;
        fc1_weights[17][83] = 16'sd-21;
        fc1_weights[17][84] = 16'sd25;
        fc1_weights[17][85] = 16'sd74;
        fc1_weights[17][86] = 16'sd59;
        fc1_weights[17][87] = 16'sd9;
        fc1_weights[17][88] = 16'sd-27;
        fc1_weights[17][89] = 16'sd54;
        fc1_weights[17][90] = 16'sd-21;
        fc1_weights[17][91] = 16'sd11;
        fc1_weights[17][92] = 16'sd1;
        fc1_weights[17][93] = 16'sd-17;
        fc1_weights[17][94] = 16'sd30;
        fc1_weights[17][95] = 16'sd55;
        fc1_weights[17][96] = 16'sd33;
        fc1_weights[17][97] = 16'sd-9;
        fc1_weights[17][98] = 16'sd89;
        fc1_weights[17][99] = 16'sd17;
        fc1_weights[17][100] = 16'sd-5;
        fc1_weights[17][101] = 16'sd-4;
        fc1_weights[17][102] = 16'sd41;
        fc1_weights[17][103] = 16'sd10;
        fc1_weights[17][104] = 16'sd-80;
        fc1_weights[17][105] = 16'sd-28;
        fc1_weights[17][106] = 16'sd6;
        fc1_weights[17][107] = 16'sd-23;
        fc1_weights[17][108] = 16'sd9;
        fc1_weights[17][109] = 16'sd11;
        fc1_weights[17][110] = 16'sd52;
        fc1_weights[17][111] = 16'sd28;
        fc1_weights[17][112] = 16'sd-34;
        fc1_weights[17][113] = 16'sd8;
        fc1_weights[17][114] = 16'sd-62;
        fc1_weights[17][115] = 16'sd-49;
        fc1_weights[17][116] = 16'sd35;
        fc1_weights[17][117] = 16'sd-11;
        fc1_weights[17][118] = 16'sd-38;
        fc1_weights[17][119] = 16'sd16;
        fc1_weights[17][120] = 16'sd48;
        fc1_weights[17][121] = 16'sd52;
        fc1_weights[17][122] = 16'sd91;
        fc1_weights[17][123] = 16'sd66;
        fc1_weights[17][124] = 16'sd89;
        fc1_weights[17][125] = 16'sd78;
        fc1_weights[17][126] = 16'sd-37;
        fc1_weights[17][127] = 16'sd-43;
        fc1_weights[17][128] = 16'sd-31;
        fc1_weights[17][129] = 16'sd9;
        fc1_weights[17][130] = 16'sd2;
        fc1_weights[17][131] = 16'sd31;
        fc1_weights[17][132] = 16'sd34;
        fc1_weights[17][133] = 16'sd18;
        fc1_weights[17][134] = 16'sd39;
        fc1_weights[17][135] = 16'sd29;
        fc1_weights[17][136] = 16'sd8;
        fc1_weights[17][137] = 16'sd-15;
        fc1_weights[17][138] = 16'sd-38;
        fc1_weights[17][139] = 16'sd10;
        fc1_weights[17][140] = 16'sd-10;
        fc1_weights[17][141] = 16'sd4;
        fc1_weights[17][142] = 16'sd63;
        fc1_weights[17][143] = 16'sd62;
        fc1_weights[17][144] = 16'sd-37;
        fc1_weights[17][145] = 16'sd-50;
        fc1_weights[17][146] = 16'sd3;
        fc1_weights[17][147] = 16'sd22;
        fc1_weights[17][148] = 16'sd-34;
        fc1_weights[17][149] = 16'sd2;
        fc1_weights[17][150] = 16'sd6;
        fc1_weights[17][151] = 16'sd-21;
        fc1_weights[17][152] = 16'sd11;
        fc1_weights[17][153] = 16'sd12;
        fc1_weights[17][154] = 16'sd45;
        fc1_weights[17][155] = 16'sd42;
        fc1_weights[17][156] = 16'sd26;
        fc1_weights[17][157] = 16'sd27;
        fc1_weights[17][158] = 16'sd41;
        fc1_weights[17][159] = 16'sd-30;
        fc1_weights[17][160] = 16'sd29;
        fc1_weights[17][161] = 16'sd39;
        fc1_weights[17][162] = 16'sd18;
        fc1_weights[17][163] = 16'sd20;
        fc1_weights[17][164] = 16'sd41;
        fc1_weights[17][165] = 16'sd48;
        fc1_weights[17][166] = 16'sd9;
        fc1_weights[17][167] = 16'sd75;
        fc1_weights[17][168] = 16'sd11;
        fc1_weights[17][169] = 16'sd47;
        fc1_weights[17][170] = 16'sd47;
        fc1_weights[17][171] = 16'sd42;
        fc1_weights[17][172] = 16'sd-27;
        fc1_weights[17][173] = 16'sd36;
        fc1_weights[17][174] = 16'sd46;
        fc1_weights[17][175] = 16'sd112;
        fc1_weights[17][176] = 16'sd90;
        fc1_weights[17][177] = 16'sd17;
        fc1_weights[17][178] = 16'sd3;
        fc1_weights[17][179] = 16'sd56;
        fc1_weights[17][180] = 16'sd45;
        fc1_weights[17][181] = 16'sd-45;
        fc1_weights[17][182] = 16'sd-53;
        fc1_weights[17][183] = 16'sd-28;
        fc1_weights[17][184] = 16'sd18;
        fc1_weights[17][185] = 16'sd-18;
        fc1_weights[17][186] = 16'sd-41;
        fc1_weights[17][187] = 16'sd-1;
        fc1_weights[17][188] = 16'sd8;
        fc1_weights[17][189] = 16'sd7;
        fc1_weights[17][190] = 16'sd6;
        fc1_weights[17][191] = 16'sd6;
        fc1_weights[17][192] = 16'sd26;
        fc1_weights[17][193] = 16'sd7;
        fc1_weights[17][194] = 16'sd11;
        fc1_weights[17][195] = 16'sd-7;
        fc1_weights[17][196] = 16'sd51;
        fc1_weights[17][197] = 16'sd-35;
        fc1_weights[17][198] = 16'sd60;
        fc1_weights[17][199] = 16'sd-4;
        fc1_weights[17][200] = 16'sd-34;
        fc1_weights[17][201] = 16'sd-3;
        fc1_weights[17][202] = 16'sd13;
        fc1_weights[17][203] = 16'sd-41;
        fc1_weights[17][204] = 16'sd-5;
        fc1_weights[17][205] = 16'sd-58;
        fc1_weights[17][206] = 16'sd-23;
        fc1_weights[17][207] = 16'sd-41;
        fc1_weights[18][0] = 16'sd43;
        fc1_weights[18][1] = 16'sd30;
        fc1_weights[18][2] = 16'sd65;
        fc1_weights[18][3] = 16'sd29;
        fc1_weights[18][4] = 16'sd9;
        fc1_weights[18][5] = 16'sd-30;
        fc1_weights[18][6] = 16'sd14;
        fc1_weights[18][7] = 16'sd14;
        fc1_weights[18][8] = 16'sd-15;
        fc1_weights[18][9] = 16'sd-51;
        fc1_weights[18][10] = 16'sd-14;
        fc1_weights[18][11] = 16'sd-55;
        fc1_weights[18][12] = 16'sd-16;
        fc1_weights[18][13] = 16'sd-9;
        fc1_weights[18][14] = 16'sd-2;
        fc1_weights[18][15] = 16'sd-19;
        fc1_weights[18][16] = 16'sd35;
        fc1_weights[18][17] = 16'sd86;
        fc1_weights[18][18] = 16'sd51;
        fc1_weights[18][19] = 16'sd24;
        fc1_weights[18][20] = 16'sd8;
        fc1_weights[18][21] = 16'sd61;
        fc1_weights[18][22] = 16'sd38;
        fc1_weights[18][23] = 16'sd44;
        fc1_weights[18][24] = 16'sd-2;
        fc1_weights[18][25] = 16'sd45;
        fc1_weights[18][26] = 16'sd15;
        fc1_weights[18][27] = 16'sd12;
        fc1_weights[18][28] = 16'sd-40;
        fc1_weights[18][29] = 16'sd22;
        fc1_weights[18][30] = 16'sd15;
        fc1_weights[18][31] = 16'sd31;
        fc1_weights[18][32] = 16'sd-14;
        fc1_weights[18][33] = 16'sd16;
        fc1_weights[18][34] = 16'sd16;
        fc1_weights[18][35] = 16'sd9;
        fc1_weights[18][36] = 16'sd8;
        fc1_weights[18][37] = 16'sd14;
        fc1_weights[18][38] = 16'sd-37;
        fc1_weights[18][39] = 16'sd-22;
        fc1_weights[18][40] = 16'sd-13;
        fc1_weights[18][41] = 16'sd-8;
        fc1_weights[18][42] = 16'sd12;
        fc1_weights[18][43] = 16'sd55;
        fc1_weights[18][44] = 16'sd-5;
        fc1_weights[18][45] = 16'sd-18;
        fc1_weights[18][46] = 16'sd-18;
        fc1_weights[18][47] = 16'sd-19;
        fc1_weights[18][48] = 16'sd0;
        fc1_weights[18][49] = 16'sd-24;
        fc1_weights[18][50] = 16'sd9;
        fc1_weights[18][51] = 16'sd-16;
        fc1_weights[18][52] = 16'sd21;
        fc1_weights[18][53] = 16'sd9;
        fc1_weights[18][54] = 16'sd-7;
        fc1_weights[18][55] = 16'sd-4;
        fc1_weights[18][56] = 16'sd-59;
        fc1_weights[18][57] = 16'sd13;
        fc1_weights[18][58] = 16'sd30;
        fc1_weights[18][59] = 16'sd27;
        fc1_weights[18][60] = 16'sd35;
        fc1_weights[18][61] = 16'sd40;
        fc1_weights[18][62] = 16'sd13;
        fc1_weights[18][63] = 16'sd1;
        fc1_weights[18][64] = 16'sd9;
        fc1_weights[18][65] = 16'sd9;
        fc1_weights[18][66] = 16'sd-26;
        fc1_weights[18][67] = 16'sd-18;
        fc1_weights[18][68] = 16'sd9;
        fc1_weights[18][69] = 16'sd-34;
        fc1_weights[18][70] = 16'sd-17;
        fc1_weights[18][71] = 16'sd-31;
        fc1_weights[18][72] = 16'sd-24;
        fc1_weights[18][73] = 16'sd-8;
        fc1_weights[18][74] = 16'sd-16;
        fc1_weights[18][75] = 16'sd13;
        fc1_weights[18][76] = 16'sd-9;
        fc1_weights[18][77] = 16'sd-26;
        fc1_weights[18][78] = 16'sd3;
        fc1_weights[18][79] = 16'sd15;
        fc1_weights[18][80] = 16'sd11;
        fc1_weights[18][81] = 16'sd12;
        fc1_weights[18][82] = 16'sd-19;
        fc1_weights[18][83] = 16'sd-35;
        fc1_weights[18][84] = 16'sd9;
        fc1_weights[18][85] = 16'sd-18;
        fc1_weights[18][86] = 16'sd-60;
        fc1_weights[18][87] = 16'sd-32;
        fc1_weights[18][88] = 16'sd7;
        fc1_weights[18][89] = 16'sd-9;
        fc1_weights[18][90] = 16'sd-32;
        fc1_weights[18][91] = 16'sd15;
        fc1_weights[18][92] = 16'sd-9;
        fc1_weights[18][93] = 16'sd-2;
        fc1_weights[18][94] = 16'sd-5;
        fc1_weights[18][95] = 16'sd16;
        fc1_weights[18][96] = 16'sd-15;
        fc1_weights[18][97] = 16'sd-7;
        fc1_weights[18][98] = 16'sd-23;
        fc1_weights[18][99] = 16'sd-35;
        fc1_weights[18][100] = 16'sd5;
        fc1_weights[18][101] = 16'sd-5;
        fc1_weights[18][102] = 16'sd-3;
        fc1_weights[18][103] = 16'sd-3;
        fc1_weights[18][104] = 16'sd-12;
        fc1_weights[18][105] = 16'sd3;
        fc1_weights[18][106] = 16'sd20;
        fc1_weights[18][107] = 16'sd-55;
        fc1_weights[18][108] = 16'sd15;
        fc1_weights[18][109] = 16'sd-14;
        fc1_weights[18][110] = 16'sd-3;
        fc1_weights[18][111] = 16'sd-39;
        fc1_weights[18][112] = 16'sd-90;
        fc1_weights[18][113] = 16'sd-123;
        fc1_weights[18][114] = 16'sd-1;
        fc1_weights[18][115] = 16'sd-6;
        fc1_weights[18][116] = 16'sd-61;
        fc1_weights[18][117] = 16'sd-69;
        fc1_weights[18][118] = 16'sd-54;
        fc1_weights[18][119] = 16'sd-32;
        fc1_weights[18][120] = 16'sd-46;
        fc1_weights[18][121] = 16'sd-29;
        fc1_weights[18][122] = 16'sd-42;
        fc1_weights[18][123] = 16'sd-70;
        fc1_weights[18][124] = 16'sd-9;
        fc1_weights[18][125] = 16'sd-9;
        fc1_weights[18][126] = 16'sd19;
        fc1_weights[18][127] = 16'sd-9;
        fc1_weights[18][128] = 16'sd19;
        fc1_weights[18][129] = 16'sd-8;
        fc1_weights[18][130] = 16'sd-39;
        fc1_weights[18][131] = 16'sd2;
        fc1_weights[18][132] = 16'sd-23;
        fc1_weights[18][133] = 16'sd-7;
        fc1_weights[18][134] = 16'sd59;
        fc1_weights[18][135] = 16'sd13;
        fc1_weights[18][136] = 16'sd54;
        fc1_weights[18][137] = 16'sd34;
        fc1_weights[18][138] = 16'sd49;
        fc1_weights[18][139] = 16'sd49;
        fc1_weights[18][140] = 16'sd96;
        fc1_weights[18][141] = 16'sd74;
        fc1_weights[18][142] = 16'sd29;
        fc1_weights[18][143] = 16'sd35;
        fc1_weights[18][144] = 16'sd47;
        fc1_weights[18][145] = 16'sd37;
        fc1_weights[18][146] = 16'sd20;
        fc1_weights[18][147] = 16'sd19;
        fc1_weights[18][148] = 16'sd-18;
        fc1_weights[18][149] = 16'sd26;
        fc1_weights[18][150] = 16'sd-13;
        fc1_weights[18][151] = 16'sd5;
        fc1_weights[18][152] = 16'sd57;
        fc1_weights[18][153] = 16'sd-9;
        fc1_weights[18][154] = 16'sd22;
        fc1_weights[18][155] = 16'sd-25;
        fc1_weights[18][156] = 16'sd55;
        fc1_weights[18][157] = 16'sd37;
        fc1_weights[18][158] = 16'sd15;
        fc1_weights[18][159] = 16'sd14;
        fc1_weights[18][160] = 16'sd49;
        fc1_weights[18][161] = 16'sd7;
        fc1_weights[18][162] = 16'sd-5;
        fc1_weights[18][163] = 16'sd16;
        fc1_weights[18][164] = 16'sd22;
        fc1_weights[18][165] = 16'sd49;
        fc1_weights[18][166] = 16'sd33;
        fc1_weights[18][167] = 16'sd-4;
        fc1_weights[18][168] = 16'sd5;
        fc1_weights[18][169] = 16'sd-12;
        fc1_weights[18][170] = 16'sd-30;
        fc1_weights[18][171] = 16'sd-23;
        fc1_weights[18][172] = 16'sd26;
        fc1_weights[18][173] = 16'sd4;
        fc1_weights[18][174] = 16'sd14;
        fc1_weights[18][175] = 16'sd8;
        fc1_weights[18][176] = 16'sd20;
        fc1_weights[18][177] = 16'sd-6;
        fc1_weights[18][178] = 16'sd20;
        fc1_weights[18][179] = 16'sd3;
        fc1_weights[18][180] = 16'sd-21;
        fc1_weights[18][181] = 16'sd4;
        fc1_weights[18][182] = 16'sd57;
        fc1_weights[18][183] = 16'sd42;
        fc1_weights[18][184] = 16'sd37;
        fc1_weights[18][185] = 16'sd9;
        fc1_weights[18][186] = 16'sd-22;
        fc1_weights[18][187] = 16'sd-22;
        fc1_weights[18][188] = 16'sd25;
        fc1_weights[18][189] = 16'sd-26;
        fc1_weights[18][190] = 16'sd-1;
        fc1_weights[18][191] = 16'sd-15;
        fc1_weights[18][192] = 16'sd5;
        fc1_weights[18][193] = 16'sd2;
        fc1_weights[18][194] = 16'sd-18;
        fc1_weights[18][195] = 16'sd1;
        fc1_weights[18][196] = 16'sd-11;
        fc1_weights[18][197] = 16'sd-35;
        fc1_weights[18][198] = 16'sd-34;
        fc1_weights[18][199] = 16'sd-22;
        fc1_weights[18][200] = 16'sd-12;
        fc1_weights[18][201] = 16'sd4;
        fc1_weights[18][202] = 16'sd-17;
        fc1_weights[18][203] = 16'sd-11;
        fc1_weights[18][204] = 16'sd-2;
        fc1_weights[18][205] = 16'sd36;
        fc1_weights[18][206] = 16'sd-2;
        fc1_weights[18][207] = 16'sd6;
        fc1_weights[19][0] = 16'sd17;
        fc1_weights[19][1] = 16'sd11;
        fc1_weights[19][2] = 16'sd6;
        fc1_weights[19][3] = 16'sd6;
        fc1_weights[19][4] = 16'sd-3;
        fc1_weights[19][5] = 16'sd5;
        fc1_weights[19][6] = 16'sd26;
        fc1_weights[19][7] = 16'sd9;
        fc1_weights[19][8] = 16'sd-6;
        fc1_weights[19][9] = 16'sd15;
        fc1_weights[19][10] = 16'sd22;
        fc1_weights[19][11] = 16'sd52;
        fc1_weights[19][12] = 16'sd-26;
        fc1_weights[19][13] = 16'sd-25;
        fc1_weights[19][14] = 16'sd6;
        fc1_weights[19][15] = 16'sd8;
        fc1_weights[19][16] = 16'sd17;
        fc1_weights[19][17] = 16'sd-29;
        fc1_weights[19][18] = 16'sd-14;
        fc1_weights[19][19] = 16'sd12;
        fc1_weights[19][20] = 16'sd56;
        fc1_weights[19][21] = 16'sd2;
        fc1_weights[19][22] = 16'sd21;
        fc1_weights[19][23] = 16'sd-20;
        fc1_weights[19][24] = 16'sd36;
        fc1_weights[19][25] = 16'sd8;
        fc1_weights[19][26] = 16'sd-15;
        fc1_weights[19][27] = 16'sd19;
        fc1_weights[19][28] = 16'sd8;
        fc1_weights[19][29] = 16'sd18;
        fc1_weights[19][30] = 16'sd12;
        fc1_weights[19][31] = 16'sd10;
        fc1_weights[19][32] = 16'sd40;
        fc1_weights[19][33] = 16'sd22;
        fc1_weights[19][34] = 16'sd-16;
        fc1_weights[19][35] = 16'sd-23;
        fc1_weights[19][36] = 16'sd45;
        fc1_weights[19][37] = 16'sd-15;
        fc1_weights[19][38] = 16'sd-31;
        fc1_weights[19][39] = 16'sd-19;
        fc1_weights[19][40] = 16'sd32;
        fc1_weights[19][41] = 16'sd-3;
        fc1_weights[19][42] = 16'sd-18;
        fc1_weights[19][43] = 16'sd36;
        fc1_weights[19][44] = 16'sd9;
        fc1_weights[19][45] = 16'sd17;
        fc1_weights[19][46] = 16'sd37;
        fc1_weights[19][47] = 16'sd28;
        fc1_weights[19][48] = 16'sd22;
        fc1_weights[19][49] = 16'sd-9;
        fc1_weights[19][50] = 16'sd4;
        fc1_weights[19][51] = 16'sd-1;
        fc1_weights[19][52] = 16'sd-31;
        fc1_weights[19][53] = 16'sd10;
        fc1_weights[19][54] = 16'sd19;
        fc1_weights[19][55] = 16'sd36;
        fc1_weights[19][56] = 16'sd-4;
        fc1_weights[19][57] = 16'sd28;
        fc1_weights[19][58] = 16'sd43;
        fc1_weights[19][59] = 16'sd25;
        fc1_weights[19][60] = 16'sd24;
        fc1_weights[19][61] = 16'sd16;
        fc1_weights[19][62] = 16'sd14;
        fc1_weights[19][63] = 16'sd10;
        fc1_weights[19][64] = 16'sd-18;
        fc1_weights[19][65] = 16'sd-4;
        fc1_weights[19][66] = 16'sd-30;
        fc1_weights[19][67] = 16'sd1;
        fc1_weights[19][68] = 16'sd19;
        fc1_weights[19][69] = 16'sd36;
        fc1_weights[19][70] = 16'sd20;
        fc1_weights[19][71] = 16'sd37;
        fc1_weights[19][72] = 16'sd39;
        fc1_weights[19][73] = 16'sd-4;
        fc1_weights[19][74] = 16'sd3;
        fc1_weights[19][75] = 16'sd-2;
        fc1_weights[19][76] = 16'sd31;
        fc1_weights[19][77] = 16'sd7;
        fc1_weights[19][78] = 16'sd-2;
        fc1_weights[19][79] = 16'sd47;
        fc1_weights[19][80] = 16'sd-10;
        fc1_weights[19][81] = 16'sd-8;
        fc1_weights[19][82] = 16'sd-18;
        fc1_weights[19][83] = 16'sd-20;
        fc1_weights[19][84] = 16'sd-2;
        fc1_weights[19][85] = 16'sd9;
        fc1_weights[19][86] = 16'sd-7;
        fc1_weights[19][87] = 16'sd-6;
        fc1_weights[19][88] = 16'sd-10;
        fc1_weights[19][89] = 16'sd7;
        fc1_weights[19][90] = 16'sd13;
        fc1_weights[19][91] = 16'sd17;
        fc1_weights[19][92] = 16'sd-8;
        fc1_weights[19][93] = 16'sd-16;
        fc1_weights[19][94] = 16'sd2;
        fc1_weights[19][95] = 16'sd12;
        fc1_weights[19][96] = 16'sd16;
        fc1_weights[19][97] = 16'sd8;
        fc1_weights[19][98] = 16'sd12;
        fc1_weights[19][99] = 16'sd-1;
        fc1_weights[19][100] = 16'sd6;
        fc1_weights[19][101] = 16'sd10;
        fc1_weights[19][102] = 16'sd23;
        fc1_weights[19][103] = 16'sd13;
        fc1_weights[19][104] = 16'sd-13;
        fc1_weights[19][105] = 16'sd-22;
        fc1_weights[19][106] = 16'sd-47;
        fc1_weights[19][107] = 16'sd-18;
        fc1_weights[19][108] = 16'sd-21;
        fc1_weights[19][109] = 16'sd-19;
        fc1_weights[19][110] = 16'sd-1;
        fc1_weights[19][111] = 16'sd-6;
        fc1_weights[19][112] = 16'sd-31;
        fc1_weights[19][113] = 16'sd-14;
        fc1_weights[19][114] = 16'sd49;
        fc1_weights[19][115] = 16'sd15;
        fc1_weights[19][116] = 16'sd86;
        fc1_weights[19][117] = 16'sd-14;
        fc1_weights[19][118] = 16'sd-38;
        fc1_weights[19][119] = 16'sd0;
        fc1_weights[19][120] = 16'sd-27;
        fc1_weights[19][121] = 16'sd0;
        fc1_weights[19][122] = 16'sd6;
        fc1_weights[19][123] = 16'sd-19;
        fc1_weights[19][124] = 16'sd-10;
        fc1_weights[19][125] = 16'sd36;
        fc1_weights[19][126] = 16'sd-8;
        fc1_weights[19][127] = 16'sd-16;
        fc1_weights[19][128] = 16'sd-34;
        fc1_weights[19][129] = 16'sd-56;
        fc1_weights[19][130] = 16'sd40;
        fc1_weights[19][131] = 16'sd17;
        fc1_weights[19][132] = 16'sd8;
        fc1_weights[19][133] = 16'sd7;
        fc1_weights[19][134] = 16'sd11;
        fc1_weights[19][135] = 16'sd-5;
        fc1_weights[19][136] = 16'sd-7;
        fc1_weights[19][137] = 16'sd1;
        fc1_weights[19][138] = 16'sd-21;
        fc1_weights[19][139] = 16'sd27;
        fc1_weights[19][140] = 16'sd25;
        fc1_weights[19][141] = 16'sd-26;
        fc1_weights[19][142] = 16'sd21;
        fc1_weights[19][143] = 16'sd4;
        fc1_weights[19][144] = 16'sd-34;
        fc1_weights[19][145] = 16'sd-34;
        fc1_weights[19][146] = 16'sd-17;
        fc1_weights[19][147] = 16'sd15;
        fc1_weights[19][148] = 16'sd-25;
        fc1_weights[19][149] = 16'sd-36;
        fc1_weights[19][150] = 16'sd-66;
        fc1_weights[19][151] = 16'sd17;
        fc1_weights[19][152] = 16'sd-28;
        fc1_weights[19][153] = 16'sd-15;
        fc1_weights[19][154] = 16'sd-20;
        fc1_weights[19][155] = 16'sd39;
        fc1_weights[19][156] = 16'sd-1;
        fc1_weights[19][157] = 16'sd-24;
        fc1_weights[19][158] = 16'sd-6;
        fc1_weights[19][159] = 16'sd7;
        fc1_weights[19][160] = 16'sd-49;
        fc1_weights[19][161] = 16'sd3;
        fc1_weights[19][162] = 16'sd-7;
        fc1_weights[19][163] = 16'sd18;
        fc1_weights[19][164] = 16'sd2;
        fc1_weights[19][165] = 16'sd-3;
        fc1_weights[19][166] = 16'sd33;
        fc1_weights[19][167] = 16'sd21;
        fc1_weights[19][168] = 16'sd-22;
        fc1_weights[19][169] = 16'sd3;
        fc1_weights[19][170] = 16'sd-8;
        fc1_weights[19][171] = 16'sd20;
        fc1_weights[19][172] = 16'sd-14;
        fc1_weights[19][173] = 16'sd-19;
        fc1_weights[19][174] = 16'sd-19;
        fc1_weights[19][175] = 16'sd36;
        fc1_weights[19][176] = 16'sd19;
        fc1_weights[19][177] = 16'sd-24;
        fc1_weights[19][178] = 16'sd-5;
        fc1_weights[19][179] = 16'sd19;
        fc1_weights[19][180] = 16'sd-1;
        fc1_weights[19][181] = 16'sd-23;
        fc1_weights[19][182] = 16'sd9;
        fc1_weights[19][183] = 16'sd-4;
        fc1_weights[19][184] = 16'sd13;
        fc1_weights[19][185] = 16'sd32;
        fc1_weights[19][186] = 16'sd-53;
        fc1_weights[19][187] = 16'sd-18;
        fc1_weights[19][188] = 16'sd20;
        fc1_weights[19][189] = 16'sd2;
        fc1_weights[19][190] = 16'sd17;
        fc1_weights[19][191] = 16'sd14;
        fc1_weights[19][192] = 16'sd-10;
        fc1_weights[19][193] = 16'sd6;
        fc1_weights[19][194] = 16'sd0;
        fc1_weights[19][195] = 16'sd-16;
        fc1_weights[19][196] = 16'sd2;
        fc1_weights[19][197] = 16'sd15;
        fc1_weights[19][198] = 16'sd19;
        fc1_weights[19][199] = 16'sd-14;
        fc1_weights[19][200] = 16'sd-27;
        fc1_weights[19][201] = 16'sd7;
        fc1_weights[19][202] = 16'sd-16;
        fc1_weights[19][203] = 16'sd-29;
        fc1_weights[19][204] = 16'sd-23;
        fc1_weights[19][205] = 16'sd17;
        fc1_weights[19][206] = 16'sd-13;
        fc1_weights[19][207] = 16'sd9;
        fc1_weights[20][0] = 16'sd7;
        fc1_weights[20][1] = 16'sd-12;
        fc1_weights[20][2] = 16'sd34;
        fc1_weights[20][3] = 16'sd19;
        fc1_weights[20][4] = 16'sd51;
        fc1_weights[20][5] = 16'sd48;
        fc1_weights[20][6] = 16'sd60;
        fc1_weights[20][7] = 16'sd4;
        fc1_weights[20][8] = 16'sd73;
        fc1_weights[20][9] = 16'sd50;
        fc1_weights[20][10] = 16'sd57;
        fc1_weights[20][11] = 16'sd51;
        fc1_weights[20][12] = 16'sd12;
        fc1_weights[20][13] = 16'sd1;
        fc1_weights[20][14] = 16'sd-15;
        fc1_weights[20][15] = 16'sd37;
        fc1_weights[20][16] = 16'sd-11;
        fc1_weights[20][17] = 16'sd-42;
        fc1_weights[20][18] = 16'sd3;
        fc1_weights[20][19] = 16'sd-5;
        fc1_weights[20][20] = 16'sd-13;
        fc1_weights[20][21] = 16'sd36;
        fc1_weights[20][22] = 16'sd48;
        fc1_weights[20][23] = 16'sd48;
        fc1_weights[20][24] = 16'sd25;
        fc1_weights[20][25] = 16'sd25;
        fc1_weights[20][26] = 16'sd40;
        fc1_weights[20][27] = 16'sd-26;
        fc1_weights[20][28] = 16'sd44;
        fc1_weights[20][29] = 16'sd-27;
        fc1_weights[20][30] = 16'sd-32;
        fc1_weights[20][31] = 16'sd5;
        fc1_weights[20][32] = 16'sd-32;
        fc1_weights[20][33] = 16'sd38;
        fc1_weights[20][34] = 16'sd-27;
        fc1_weights[20][35] = 16'sd-67;
        fc1_weights[20][36] = 16'sd17;
        fc1_weights[20][37] = 16'sd28;
        fc1_weights[20][38] = 16'sd-36;
        fc1_weights[20][39] = 16'sd-25;
        fc1_weights[20][40] = 16'sd-11;
        fc1_weights[20][41] = 16'sd-18;
        fc1_weights[20][42] = 16'sd41;
        fc1_weights[20][43] = 16'sd23;
        fc1_weights[20][44] = 16'sd8;
        fc1_weights[20][45] = 16'sd8;
        fc1_weights[20][46] = 16'sd-3;
        fc1_weights[20][47] = 16'sd18;
        fc1_weights[20][48] = 16'sd-22;
        fc1_weights[20][49] = 16'sd-20;
        fc1_weights[20][50] = 16'sd-21;
        fc1_weights[20][51] = 16'sd7;
        fc1_weights[20][52] = 16'sd-26;
        fc1_weights[20][53] = 16'sd-23;
        fc1_weights[20][54] = 16'sd10;
        fc1_weights[20][55] = 16'sd-34;
        fc1_weights[20][56] = 16'sd-18;
        fc1_weights[20][57] = 16'sd-35;
        fc1_weights[20][58] = 16'sd-62;
        fc1_weights[20][59] = 16'sd-23;
        fc1_weights[20][60] = 16'sd-72;
        fc1_weights[20][61] = 16'sd-92;
        fc1_weights[20][62] = 16'sd-47;
        fc1_weights[20][63] = 16'sd23;
        fc1_weights[20][64] = 16'sd-79;
        fc1_weights[20][65] = 16'sd-3;
        fc1_weights[20][66] = 16'sd49;
        fc1_weights[20][67] = 16'sd9;
        fc1_weights[20][68] = 16'sd62;
        fc1_weights[20][69] = 16'sd-33;
        fc1_weights[20][70] = 16'sd-43;
        fc1_weights[20][71] = 16'sd-58;
        fc1_weights[20][72] = 16'sd10;
        fc1_weights[20][73] = 16'sd20;
        fc1_weights[20][74] = 16'sd-9;
        fc1_weights[20][75] = 16'sd45;
        fc1_weights[20][76] = 16'sd-17;
        fc1_weights[20][77] = 16'sd-39;
        fc1_weights[20][78] = 16'sd-89;
        fc1_weights[20][79] = 16'sd29;
        fc1_weights[20][80] = 16'sd0;
        fc1_weights[20][81] = 16'sd-19;
        fc1_weights[20][82] = 16'sd2;
        fc1_weights[20][83] = 16'sd-95;
        fc1_weights[20][84] = 16'sd-28;
        fc1_weights[20][85] = 16'sd8;
        fc1_weights[20][86] = 16'sd-3;
        fc1_weights[20][87] = 16'sd-62;
        fc1_weights[20][88] = 16'sd-35;
        fc1_weights[20][89] = 16'sd64;
        fc1_weights[20][90] = 16'sd-36;
        fc1_weights[20][91] = 16'sd-9;
        fc1_weights[20][92] = 16'sd-39;
        fc1_weights[20][93] = 16'sd-32;
        fc1_weights[20][94] = 16'sd0;
        fc1_weights[20][95] = 16'sd-28;
        fc1_weights[20][96] = 16'sd9;
        fc1_weights[20][97] = 16'sd8;
        fc1_weights[20][98] = 16'sd63;
        fc1_weights[20][99] = 16'sd88;
        fc1_weights[20][100] = 16'sd2;
        fc1_weights[20][101] = 16'sd45;
        fc1_weights[20][102] = 16'sd46;
        fc1_weights[20][103] = 16'sd12;
        fc1_weights[20][104] = 16'sd-56;
        fc1_weights[20][105] = 16'sd10;
        fc1_weights[20][106] = 16'sd-6;
        fc1_weights[20][107] = 16'sd-19;
        fc1_weights[20][108] = 16'sd-12;
        fc1_weights[20][109] = 16'sd-39;
        fc1_weights[20][110] = 16'sd4;
        fc1_weights[20][111] = 16'sd-5;
        fc1_weights[20][112] = 16'sd-35;
        fc1_weights[20][113] = 16'sd-19;
        fc1_weights[20][114] = 16'sd-37;
        fc1_weights[20][115] = 16'sd-17;
        fc1_weights[20][116] = 16'sd-57;
        fc1_weights[20][117] = 16'sd11;
        fc1_weights[20][118] = 16'sd-14;
        fc1_weights[20][119] = 16'sd34;
        fc1_weights[20][120] = 16'sd41;
        fc1_weights[20][121] = 16'sd18;
        fc1_weights[20][122] = 16'sd35;
        fc1_weights[20][123] = 16'sd15;
        fc1_weights[20][124] = 16'sd66;
        fc1_weights[20][125] = 16'sd-2;
        fc1_weights[20][126] = 16'sd19;
        fc1_weights[20][127] = 16'sd-21;
        fc1_weights[20][128] = 16'sd-29;
        fc1_weights[20][129] = 16'sd-2;
        fc1_weights[20][130] = 16'sd-27;
        fc1_weights[20][131] = 16'sd5;
        fc1_weights[20][132] = 16'sd4;
        fc1_weights[20][133] = 16'sd11;
        fc1_weights[20][134] = 16'sd37;
        fc1_weights[20][135] = 16'sd42;
        fc1_weights[20][136] = 16'sd64;
        fc1_weights[20][137] = 16'sd29;
        fc1_weights[20][138] = 16'sd-21;
        fc1_weights[20][139] = 16'sd61;
        fc1_weights[20][140] = 16'sd15;
        fc1_weights[20][141] = 16'sd19;
        fc1_weights[20][142] = 16'sd27;
        fc1_weights[20][143] = 16'sd43;
        fc1_weights[20][144] = 16'sd-58;
        fc1_weights[20][145] = 16'sd-5;
        fc1_weights[20][146] = 16'sd4;
        fc1_weights[20][147] = 16'sd-5;
        fc1_weights[20][148] = 16'sd21;
        fc1_weights[20][149] = 16'sd38;
        fc1_weights[20][150] = 16'sd3;
        fc1_weights[20][151] = 16'sd-18;
        fc1_weights[20][152] = 16'sd17;
        fc1_weights[20][153] = 16'sd2;
        fc1_weights[20][154] = 16'sd35;
        fc1_weights[20][155] = 16'sd7;
        fc1_weights[20][156] = 16'sd25;
        fc1_weights[20][157] = 16'sd0;
        fc1_weights[20][158] = 16'sd65;
        fc1_weights[20][159] = 16'sd13;
        fc1_weights[20][160] = 16'sd45;
        fc1_weights[20][161] = 16'sd1;
        fc1_weights[20][162] = 16'sd-17;
        fc1_weights[20][163] = 16'sd2;
        fc1_weights[20][164] = 16'sd2;
        fc1_weights[20][165] = 16'sd17;
        fc1_weights[20][166] = 16'sd-24;
        fc1_weights[20][167] = 16'sd-3;
        fc1_weights[20][168] = 16'sd17;
        fc1_weights[20][169] = 16'sd20;
        fc1_weights[20][170] = 16'sd54;
        fc1_weights[20][171] = 16'sd38;
        fc1_weights[20][172] = 16'sd34;
        fc1_weights[20][173] = 16'sd47;
        fc1_weights[20][174] = 16'sd76;
        fc1_weights[20][175] = 16'sd16;
        fc1_weights[20][176] = 16'sd39;
        fc1_weights[20][177] = 16'sd23;
        fc1_weights[20][178] = 16'sd35;
        fc1_weights[20][179] = 16'sd15;
        fc1_weights[20][180] = 16'sd39;
        fc1_weights[20][181] = 16'sd0;
        fc1_weights[20][182] = 16'sd-5;
        fc1_weights[20][183] = 16'sd14;
        fc1_weights[20][184] = 16'sd11;
        fc1_weights[20][185] = 16'sd-27;
        fc1_weights[20][186] = 16'sd-40;
        fc1_weights[20][187] = 16'sd-45;
        fc1_weights[20][188] = 16'sd-11;
        fc1_weights[20][189] = 16'sd-31;
        fc1_weights[20][190] = 16'sd16;
        fc1_weights[20][191] = 16'sd-43;
        fc1_weights[20][192] = 16'sd4;
        fc1_weights[20][193] = 16'sd33;
        fc1_weights[20][194] = 16'sd-27;
        fc1_weights[20][195] = 16'sd10;
        fc1_weights[20][196] = 16'sd18;
        fc1_weights[20][197] = 16'sd-13;
        fc1_weights[20][198] = 16'sd44;
        fc1_weights[20][199] = 16'sd4;
        fc1_weights[20][200] = 16'sd5;
        fc1_weights[20][201] = 16'sd32;
        fc1_weights[20][202] = 16'sd-24;
        fc1_weights[20][203] = 16'sd-3;
        fc1_weights[20][204] = 16'sd7;
        fc1_weights[20][205] = 16'sd-23;
        fc1_weights[20][206] = 16'sd21;
        fc1_weights[20][207] = 16'sd27;
        fc1_weights[21][0] = 16'sd14;
        fc1_weights[21][1] = 16'sd9;
        fc1_weights[21][2] = 16'sd-2;
        fc1_weights[21][3] = 16'sd8;
        fc1_weights[21][4] = 16'sd3;
        fc1_weights[21][5] = 16'sd24;
        fc1_weights[21][6] = 16'sd3;
        fc1_weights[21][7] = 16'sd9;
        fc1_weights[21][8] = 16'sd13;
        fc1_weights[21][9] = 16'sd7;
        fc1_weights[21][10] = 16'sd24;
        fc1_weights[21][11] = 16'sd5;
        fc1_weights[21][12] = 16'sd-15;
        fc1_weights[21][13] = 16'sd-18;
        fc1_weights[21][14] = 16'sd13;
        fc1_weights[21][15] = 16'sd20;
        fc1_weights[21][16] = 16'sd21;
        fc1_weights[21][17] = 16'sd6;
        fc1_weights[21][18] = 16'sd-2;
        fc1_weights[21][19] = 16'sd18;
        fc1_weights[21][20] = 16'sd32;
        fc1_weights[21][21] = 16'sd8;
        fc1_weights[21][22] = 16'sd-3;
        fc1_weights[21][23] = 16'sd6;
        fc1_weights[21][24] = 16'sd11;
        fc1_weights[21][25] = 16'sd24;
        fc1_weights[21][26] = 16'sd-12;
        fc1_weights[21][27] = 16'sd15;
        fc1_weights[21][28] = 16'sd-10;
        fc1_weights[21][29] = 16'sd3;
        fc1_weights[21][30] = 16'sd2;
        fc1_weights[21][31] = 16'sd25;
        fc1_weights[21][32] = 16'sd42;
        fc1_weights[21][33] = 16'sd33;
        fc1_weights[21][34] = 16'sd15;
        fc1_weights[21][35] = 16'sd24;
        fc1_weights[21][36] = 16'sd22;
        fc1_weights[21][37] = 16'sd6;
        fc1_weights[21][38] = 16'sd-4;
        fc1_weights[21][39] = 16'sd15;
        fc1_weights[21][40] = 16'sd22;
        fc1_weights[21][41] = 16'sd29;
        fc1_weights[21][42] = 16'sd37;
        fc1_weights[21][43] = 16'sd44;
        fc1_weights[21][44] = 16'sd29;
        fc1_weights[21][45] = 16'sd39;
        fc1_weights[21][46] = 16'sd14;
        fc1_weights[21][47] = 16'sd18;
        fc1_weights[21][48] = 16'sd1;
        fc1_weights[21][49] = 16'sd28;
        fc1_weights[21][50] = 16'sd-17;
        fc1_weights[21][51] = 16'sd11;
        fc1_weights[21][52] = 16'sd-40;
        fc1_weights[21][53] = 16'sd-12;
        fc1_weights[21][54] = 16'sd2;
        fc1_weights[21][55] = 16'sd-10;
        fc1_weights[21][56] = 16'sd12;
        fc1_weights[21][57] = 16'sd-1;
        fc1_weights[21][58] = 16'sd3;
        fc1_weights[21][59] = 16'sd1;
        fc1_weights[21][60] = 16'sd-20;
        fc1_weights[21][61] = 16'sd18;
        fc1_weights[21][62] = 16'sd19;
        fc1_weights[21][63] = 16'sd11;
        fc1_weights[21][64] = 16'sd13;
        fc1_weights[21][65] = 16'sd2;
        fc1_weights[21][66] = 16'sd8;
        fc1_weights[21][67] = 16'sd4;
        fc1_weights[21][68] = 16'sd20;
        fc1_weights[21][69] = 16'sd42;
        fc1_weights[21][70] = 16'sd31;
        fc1_weights[21][71] = 16'sd-1;
        fc1_weights[21][72] = 16'sd18;
        fc1_weights[21][73] = 16'sd14;
        fc1_weights[21][74] = 16'sd3;
        fc1_weights[21][75] = 16'sd16;
        fc1_weights[21][76] = 16'sd-3;
        fc1_weights[21][77] = 16'sd12;
        fc1_weights[21][78] = 16'sd-36;
        fc1_weights[21][79] = 16'sd-52;
        fc1_weights[21][80] = 16'sd-2;
        fc1_weights[21][81] = 16'sd-6;
        fc1_weights[21][82] = 16'sd31;
        fc1_weights[21][83] = 16'sd-17;
        fc1_weights[21][84] = 16'sd-14;
        fc1_weights[21][85] = 16'sd14;
        fc1_weights[21][86] = 16'sd-21;
        fc1_weights[21][87] = 16'sd-16;
        fc1_weights[21][88] = 16'sd-3;
        fc1_weights[21][89] = 16'sd2;
        fc1_weights[21][90] = 16'sd-24;
        fc1_weights[21][91] = 16'sd-29;
        fc1_weights[21][92] = 16'sd-36;
        fc1_weights[21][93] = 16'sd7;
        fc1_weights[21][94] = 16'sd23;
        fc1_weights[21][95] = 16'sd7;
        fc1_weights[21][96] = 16'sd7;
        fc1_weights[21][97] = 16'sd-8;
        fc1_weights[21][98] = 16'sd-1;
        fc1_weights[21][99] = 16'sd6;
        fc1_weights[21][100] = 16'sd-1;
        fc1_weights[21][101] = 16'sd28;
        fc1_weights[21][102] = 16'sd4;
        fc1_weights[21][103] = 16'sd-17;
        fc1_weights[21][104] = 16'sd-26;
        fc1_weights[21][105] = 16'sd17;
        fc1_weights[21][106] = 16'sd-16;
        fc1_weights[21][107] = 16'sd24;
        fc1_weights[21][108] = 16'sd19;
        fc1_weights[21][109] = 16'sd18;
        fc1_weights[21][110] = 16'sd32;
        fc1_weights[21][111] = 16'sd12;
        fc1_weights[21][112] = 16'sd22;
        fc1_weights[21][113] = 16'sd38;
        fc1_weights[21][114] = 16'sd-15;
        fc1_weights[21][115] = 16'sd-24;
        fc1_weights[21][116] = 16'sd-22;
        fc1_weights[21][117] = 16'sd19;
        fc1_weights[21][118] = 16'sd22;
        fc1_weights[21][119] = 16'sd0;
        fc1_weights[21][120] = 16'sd-14;
        fc1_weights[21][121] = 16'sd-7;
        fc1_weights[21][122] = 16'sd-2;
        fc1_weights[21][123] = 16'sd7;
        fc1_weights[21][124] = 16'sd11;
        fc1_weights[21][125] = 16'sd6;
        fc1_weights[21][126] = 16'sd11;
        fc1_weights[21][127] = 16'sd2;
        fc1_weights[21][128] = 16'sd2;
        fc1_weights[21][129] = 16'sd-12;
        fc1_weights[21][130] = 16'sd23;
        fc1_weights[21][131] = 16'sd38;
        fc1_weights[21][132] = 16'sd33;
        fc1_weights[21][133] = 16'sd11;
        fc1_weights[21][134] = 16'sd15;
        fc1_weights[21][135] = 16'sd25;
        fc1_weights[21][136] = 16'sd-9;
        fc1_weights[21][137] = 16'sd36;
        fc1_weights[21][138] = 16'sd43;
        fc1_weights[21][139] = 16'sd38;
        fc1_weights[21][140] = 16'sd36;
        fc1_weights[21][141] = 16'sd13;
        fc1_weights[21][142] = 16'sd20;
        fc1_weights[21][143] = 16'sd68;
        fc1_weights[21][144] = 16'sd34;
        fc1_weights[21][145] = 16'sd-3;
        fc1_weights[21][146] = 16'sd-9;
        fc1_weights[21][147] = 16'sd-18;
        fc1_weights[21][148] = 16'sd-25;
        fc1_weights[21][149] = 16'sd-5;
        fc1_weights[21][150] = 16'sd14;
        fc1_weights[21][151] = 16'sd10;
        fc1_weights[21][152] = 16'sd-4;
        fc1_weights[21][153] = 16'sd-4;
        fc1_weights[21][154] = 16'sd-24;
        fc1_weights[21][155] = 16'sd-2;
        fc1_weights[21][156] = 16'sd15;
        fc1_weights[21][157] = 16'sd-11;
        fc1_weights[21][158] = 16'sd-16;
        fc1_weights[21][159] = 16'sd36;
        fc1_weights[21][160] = 16'sd31;
        fc1_weights[21][161] = 16'sd7;
        fc1_weights[21][162] = 16'sd12;
        fc1_weights[21][163] = 16'sd-12;
        fc1_weights[21][164] = 16'sd30;
        fc1_weights[21][165] = 16'sd26;
        fc1_weights[21][166] = 16'sd-1;
        fc1_weights[21][167] = 16'sd7;
        fc1_weights[21][168] = 16'sd20;
        fc1_weights[21][169] = 16'sd31;
        fc1_weights[21][170] = 16'sd23;
        fc1_weights[21][171] = 16'sd23;
        fc1_weights[21][172] = 16'sd17;
        fc1_weights[21][173] = 16'sd3;
        fc1_weights[21][174] = 16'sd-21;
        fc1_weights[21][175] = 16'sd7;
        fc1_weights[21][176] = 16'sd11;
        fc1_weights[21][177] = 16'sd10;
        fc1_weights[21][178] = 16'sd2;
        fc1_weights[21][179] = 16'sd6;
        fc1_weights[21][180] = 16'sd-12;
        fc1_weights[21][181] = 16'sd-3;
        fc1_weights[21][182] = 16'sd18;
        fc1_weights[21][183] = 16'sd-7;
        fc1_weights[21][184] = 16'sd18;
        fc1_weights[21][185] = 16'sd34;
        fc1_weights[21][186] = 16'sd30;
        fc1_weights[21][187] = 16'sd41;
        fc1_weights[21][188] = 16'sd30;
        fc1_weights[21][189] = 16'sd20;
        fc1_weights[21][190] = 16'sd16;
        fc1_weights[21][191] = 16'sd1;
        fc1_weights[21][192] = 16'sd28;
        fc1_weights[21][193] = 16'sd34;
        fc1_weights[21][194] = 16'sd8;
        fc1_weights[21][195] = 16'sd10;
        fc1_weights[21][196] = 16'sd10;
        fc1_weights[21][197] = 16'sd20;
        fc1_weights[21][198] = 16'sd25;
        fc1_weights[21][199] = 16'sd-18;
        fc1_weights[21][200] = 16'sd10;
        fc1_weights[21][201] = 16'sd4;
        fc1_weights[21][202] = 16'sd-11;
        fc1_weights[21][203] = 16'sd-6;
        fc1_weights[21][204] = 16'sd-6;
        fc1_weights[21][205] = 16'sd-11;
        fc1_weights[21][206] = 16'sd-7;
        fc1_weights[21][207] = 16'sd5;
        fc1_weights[22][0] = 16'sd0;
        fc1_weights[22][1] = 16'sd28;
        fc1_weights[22][2] = 16'sd35;
        fc1_weights[22][3] = 16'sd18;
        fc1_weights[22][4] = 16'sd-23;
        fc1_weights[22][5] = 16'sd22;
        fc1_weights[22][6] = 16'sd25;
        fc1_weights[22][7] = 16'sd52;
        fc1_weights[22][8] = 16'sd23;
        fc1_weights[22][9] = 16'sd-10;
        fc1_weights[22][10] = 16'sd26;
        fc1_weights[22][11] = 16'sd-2;
        fc1_weights[22][12] = 16'sd40;
        fc1_weights[22][13] = 16'sd31;
        fc1_weights[22][14] = 16'sd-26;
        fc1_weights[22][15] = 16'sd-2;
        fc1_weights[22][16] = 16'sd-2;
        fc1_weights[22][17] = 16'sd-14;
        fc1_weights[22][18] = 16'sd-20;
        fc1_weights[22][19] = 16'sd-23;
        fc1_weights[22][20] = 16'sd-28;
        fc1_weights[22][21] = 16'sd-25;
        fc1_weights[22][22] = 16'sd16;
        fc1_weights[22][23] = 16'sd2;
        fc1_weights[22][24] = 16'sd7;
        fc1_weights[22][25] = 16'sd44;
        fc1_weights[22][26] = 16'sd-5;
        fc1_weights[22][27] = 16'sd-12;
        fc1_weights[22][28] = 16'sd13;
        fc1_weights[22][29] = 16'sd14;
        fc1_weights[22][30] = 16'sd-11;
        fc1_weights[22][31] = 16'sd62;
        fc1_weights[22][32] = 16'sd10;
        fc1_weights[22][33] = 16'sd45;
        fc1_weights[22][34] = 16'sd44;
        fc1_weights[22][35] = 16'sd-10;
        fc1_weights[22][36] = 16'sd3;
        fc1_weights[22][37] = 16'sd29;
        fc1_weights[22][38] = 16'sd-22;
        fc1_weights[22][39] = 16'sd-55;
        fc1_weights[22][40] = 16'sd17;
        fc1_weights[22][41] = 16'sd-79;
        fc1_weights[22][42] = 16'sd-7;
        fc1_weights[22][43] = 16'sd-47;
        fc1_weights[22][44] = 16'sd-12;
        fc1_weights[22][45] = 16'sd1;
        fc1_weights[22][46] = 16'sd-7;
        fc1_weights[22][47] = 16'sd-4;
        fc1_weights[22][48] = 16'sd2;
        fc1_weights[22][49] = 16'sd30;
        fc1_weights[22][50] = 16'sd4;
        fc1_weights[22][51] = 16'sd-19;
        fc1_weights[22][52] = 16'sd23;
        fc1_weights[22][53] = 16'sd-34;
        fc1_weights[22][54] = 16'sd-19;
        fc1_weights[22][55] = 16'sd-37;
        fc1_weights[22][56] = 16'sd-28;
        fc1_weights[22][57] = 16'sd-23;
        fc1_weights[22][58] = 16'sd-45;
        fc1_weights[22][59] = 16'sd-27;
        fc1_weights[22][60] = 16'sd12;
        fc1_weights[22][61] = 16'sd12;
        fc1_weights[22][62] = 16'sd-8;
        fc1_weights[22][63] = 16'sd14;
        fc1_weights[22][64] = 16'sd-19;
        fc1_weights[22][65] = 16'sd-29;
        fc1_weights[22][66] = 16'sd56;
        fc1_weights[22][67] = 16'sd-1;
        fc1_weights[22][68] = 16'sd-73;
        fc1_weights[22][69] = 16'sd3;
        fc1_weights[22][70] = 16'sd31;
        fc1_weights[22][71] = 16'sd21;
        fc1_weights[22][72] = 16'sd35;
        fc1_weights[22][73] = 16'sd21;
        fc1_weights[22][74] = 16'sd49;
        fc1_weights[22][75] = 16'sd29;
        fc1_weights[22][76] = 16'sd5;
        fc1_weights[22][77] = 16'sd9;
        fc1_weights[22][78] = 16'sd7;
        fc1_weights[22][79] = 16'sd71;
        fc1_weights[22][80] = 16'sd-9;
        fc1_weights[22][81] = 16'sd-2;
        fc1_weights[22][82] = 16'sd-40;
        fc1_weights[22][83] = 16'sd58;
        fc1_weights[22][84] = 16'sd8;
        fc1_weights[22][85] = 16'sd-9;
        fc1_weights[22][86] = 16'sd-10;
        fc1_weights[22][87] = 16'sd27;
        fc1_weights[22][88] = 16'sd33;
        fc1_weights[22][89] = 16'sd-9;
        fc1_weights[22][90] = 16'sd-2;
        fc1_weights[22][91] = 16'sd-17;
        fc1_weights[22][92] = 16'sd-35;
        fc1_weights[22][93] = 16'sd-4;
        fc1_weights[22][94] = 16'sd-67;
        fc1_weights[22][95] = 16'sd-27;
        fc1_weights[22][96] = 16'sd-30;
        fc1_weights[22][97] = 16'sd12;
        fc1_weights[22][98] = 16'sd25;
        fc1_weights[22][99] = 16'sd-19;
        fc1_weights[22][100] = 16'sd10;
        fc1_weights[22][101] = 16'sd-1;
        fc1_weights[22][102] = 16'sd-5;
        fc1_weights[22][103] = 16'sd-8;
        fc1_weights[22][104] = 16'sd20;
        fc1_weights[22][105] = 16'sd-19;
        fc1_weights[22][106] = 16'sd15;
        fc1_weights[22][107] = 16'sd-14;
        fc1_weights[22][108] = 16'sd25;
        fc1_weights[22][109] = 16'sd19;
        fc1_weights[22][110] = 16'sd5;
        fc1_weights[22][111] = 16'sd4;
        fc1_weights[22][112] = 16'sd53;
        fc1_weights[22][113] = 16'sd44;
        fc1_weights[22][114] = 16'sd31;
        fc1_weights[22][115] = 16'sd15;
        fc1_weights[22][116] = 16'sd-23;
        fc1_weights[22][117] = 16'sd-40;
        fc1_weights[22][118] = 16'sd-44;
        fc1_weights[22][119] = 16'sd24;
        fc1_weights[22][120] = 16'sd3;
        fc1_weights[22][121] = 16'sd20;
        fc1_weights[22][122] = 16'sd-7;
        fc1_weights[22][123] = 16'sd-17;
        fc1_weights[22][124] = 16'sd12;
        fc1_weights[22][125] = 16'sd-17;
        fc1_weights[22][126] = 16'sd-39;
        fc1_weights[22][127] = 16'sd-31;
        fc1_weights[22][128] = 16'sd-14;
        fc1_weights[22][129] = 16'sd-4;
        fc1_weights[22][130] = 16'sd-7;
        fc1_weights[22][131] = 16'sd16;
        fc1_weights[22][132] = 16'sd72;
        fc1_weights[22][133] = 16'sd31;
        fc1_weights[22][134] = 16'sd26;
        fc1_weights[22][135] = 16'sd6;
        fc1_weights[22][136] = 16'sd1;
        fc1_weights[22][137] = 16'sd44;
        fc1_weights[22][138] = 16'sd-18;
        fc1_weights[22][139] = 16'sd-4;
        fc1_weights[22][140] = 16'sd-6;
        fc1_weights[22][141] = 16'sd11;
        fc1_weights[22][142] = 16'sd-15;
        fc1_weights[22][143] = 16'sd-26;
        fc1_weights[22][144] = 16'sd35;
        fc1_weights[22][145] = 16'sd15;
        fc1_weights[22][146] = 16'sd15;
        fc1_weights[22][147] = 16'sd14;
        fc1_weights[22][148] = 16'sd37;
        fc1_weights[22][149] = 16'sd-17;
        fc1_weights[22][150] = 16'sd26;
        fc1_weights[22][151] = 16'sd11;
        fc1_weights[22][152] = 16'sd-15;
        fc1_weights[22][153] = 16'sd-33;
        fc1_weights[22][154] = 16'sd9;
        fc1_weights[22][155] = 16'sd-15;
        fc1_weights[22][156] = 16'sd20;
        fc1_weights[22][157] = 16'sd14;
        fc1_weights[22][158] = 16'sd-1;
        fc1_weights[22][159] = 16'sd25;
        fc1_weights[22][160] = 16'sd66;
        fc1_weights[22][161] = 16'sd25;
        fc1_weights[22][162] = 16'sd-4;
        fc1_weights[22][163] = 16'sd-16;
        fc1_weights[22][164] = 16'sd-40;
        fc1_weights[22][165] = 16'sd9;
        fc1_weights[22][166] = 16'sd27;
        fc1_weights[22][167] = 16'sd-2;
        fc1_weights[22][168] = 16'sd-6;
        fc1_weights[22][169] = 16'sd-22;
        fc1_weights[22][170] = 16'sd-21;
        fc1_weights[22][171] = 16'sd3;
        fc1_weights[22][172] = 16'sd-60;
        fc1_weights[22][173] = 16'sd-6;
        fc1_weights[22][174] = 16'sd40;
        fc1_weights[22][175] = 16'sd-4;
        fc1_weights[22][176] = 16'sd-16;
        fc1_weights[22][177] = 16'sd50;
        fc1_weights[22][178] = 16'sd-4;
        fc1_weights[22][179] = 16'sd-16;
        fc1_weights[22][180] = 16'sd15;
        fc1_weights[22][181] = 16'sd-6;
        fc1_weights[22][182] = 16'sd9;
        fc1_weights[22][183] = 16'sd-36;
        fc1_weights[22][184] = 16'sd-16;
        fc1_weights[22][185] = 16'sd-1;
        fc1_weights[22][186] = 16'sd-57;
        fc1_weights[22][187] = 16'sd-76;
        fc1_weights[22][188] = 16'sd-13;
        fc1_weights[22][189] = 16'sd-49;
        fc1_weights[22][190] = 16'sd12;
        fc1_weights[22][191] = 16'sd17;
        fc1_weights[22][192] = 16'sd9;
        fc1_weights[22][193] = 16'sd-12;
        fc1_weights[22][194] = 16'sd29;
        fc1_weights[22][195] = 16'sd-40;
        fc1_weights[22][196] = 16'sd-35;
        fc1_weights[22][197] = 16'sd-39;
        fc1_weights[22][198] = 16'sd11;
        fc1_weights[22][199] = 16'sd-29;
        fc1_weights[22][200] = 16'sd-14;
        fc1_weights[22][201] = 16'sd0;
        fc1_weights[22][202] = 16'sd25;
        fc1_weights[22][203] = 16'sd-9;
        fc1_weights[22][204] = 16'sd-44;
        fc1_weights[22][205] = 16'sd-9;
        fc1_weights[22][206] = 16'sd50;
        fc1_weights[22][207] = 16'sd10;
        fc1_weights[23][0] = 16'sd-55;
        fc1_weights[23][1] = 16'sd6;
        fc1_weights[23][2] = 16'sd-31;
        fc1_weights[23][3] = 16'sd2;
        fc1_weights[23][4] = 16'sd-23;
        fc1_weights[23][5] = 16'sd0;
        fc1_weights[23][6] = 16'sd27;
        fc1_weights[23][7] = 16'sd41;
        fc1_weights[23][8] = 16'sd-80;
        fc1_weights[23][9] = 16'sd-93;
        fc1_weights[23][10] = 16'sd-82;
        fc1_weights[23][11] = 16'sd-31;
        fc1_weights[23][12] = 16'sd52;
        fc1_weights[23][13] = 16'sd95;
        fc1_weights[23][14] = 16'sd79;
        fc1_weights[23][15] = 16'sd22;
        fc1_weights[23][16] = 16'sd48;
        fc1_weights[23][17] = 16'sd38;
        fc1_weights[23][18] = 16'sd30;
        fc1_weights[23][19] = 16'sd21;
        fc1_weights[23][20] = 16'sd8;
        fc1_weights[23][21] = 16'sd5;
        fc1_weights[23][22] = 16'sd21;
        fc1_weights[23][23] = 16'sd25;
        fc1_weights[23][24] = 16'sd-5;
        fc1_weights[23][25] = 16'sd-6;
        fc1_weights[23][26] = 16'sd-27;
        fc1_weights[23][27] = 16'sd-44;
        fc1_weights[23][28] = 16'sd-17;
        fc1_weights[23][29] = 16'sd35;
        fc1_weights[23][30] = 16'sd16;
        fc1_weights[23][31] = 16'sd-11;
        fc1_weights[23][32] = 16'sd-7;
        fc1_weights[23][33] = 16'sd-29;
        fc1_weights[23][34] = 16'sd-8;
        fc1_weights[23][35] = 16'sd-7;
        fc1_weights[23][36] = 16'sd-24;
        fc1_weights[23][37] = 16'sd-15;
        fc1_weights[23][38] = 16'sd14;
        fc1_weights[23][39] = 16'sd54;
        fc1_weights[23][40] = 16'sd22;
        fc1_weights[23][41] = 16'sd10;
        fc1_weights[23][42] = 16'sd2;
        fc1_weights[23][43] = 16'sd-36;
        fc1_weights[23][44] = 16'sd-18;
        fc1_weights[23][45] = 16'sd-25;
        fc1_weights[23][46] = 16'sd25;
        fc1_weights[23][47] = 16'sd25;
        fc1_weights[23][48] = 16'sd-31;
        fc1_weights[23][49] = 16'sd-18;
        fc1_weights[23][50] = 16'sd-31;
        fc1_weights[23][51] = 16'sd-48;
        fc1_weights[23][52] = 16'sd-31;
        fc1_weights[23][53] = 16'sd-19;
        fc1_weights[23][54] = 16'sd-52;
        fc1_weights[23][55] = 16'sd27;
        fc1_weights[23][56] = 16'sd9;
        fc1_weights[23][57] = 16'sd-12;
        fc1_weights[23][58] = 16'sd-5;
        fc1_weights[23][59] = 16'sd15;
        fc1_weights[23][60] = 16'sd9;
        fc1_weights[23][61] = 16'sd-19;
        fc1_weights[23][62] = 16'sd-53;
        fc1_weights[23][63] = 16'sd-7;
        fc1_weights[23][64] = 16'sd78;
        fc1_weights[23][65] = 16'sd18;
        fc1_weights[23][66] = 16'sd91;
        fc1_weights[23][67] = 16'sd11;
        fc1_weights[23][68] = 16'sd-85;
        fc1_weights[23][69] = 16'sd7;
        fc1_weights[23][70] = 16'sd1;
        fc1_weights[23][71] = 16'sd30;
        fc1_weights[23][72] = 16'sd48;
        fc1_weights[23][73] = 16'sd50;
        fc1_weights[23][74] = 16'sd14;
        fc1_weights[23][75] = 16'sd-32;
        fc1_weights[23][76] = 16'sd-56;
        fc1_weights[23][77] = 16'sd1;
        fc1_weights[23][78] = 16'sd-23;
        fc1_weights[23][79] = 16'sd-3;
        fc1_weights[23][80] = 16'sd-29;
        fc1_weights[23][81] = 16'sd8;
        fc1_weights[23][82] = 16'sd-47;
        fc1_weights[23][83] = 16'sd46;
        fc1_weights[23][84] = 16'sd16;
        fc1_weights[23][85] = 16'sd27;
        fc1_weights[23][86] = 16'sd63;
        fc1_weights[23][87] = 16'sd-4;
        fc1_weights[23][88] = 16'sd-19;
        fc1_weights[23][89] = 16'sd-60;
        fc1_weights[23][90] = 16'sd-40;
        fc1_weights[23][91] = 16'sd14;
        fc1_weights[23][92] = 16'sd16;
        fc1_weights[23][93] = 16'sd21;
        fc1_weights[23][94] = 16'sd-44;
        fc1_weights[23][95] = 16'sd31;
        fc1_weights[23][96] = 16'sd-23;
        fc1_weights[23][97] = 16'sd-14;
        fc1_weights[23][98] = 16'sd10;
        fc1_weights[23][99] = 16'sd-18;
        fc1_weights[23][100] = 16'sd4;
        fc1_weights[23][101] = 16'sd-10;
        fc1_weights[23][102] = 16'sd-44;
        fc1_weights[23][103] = 16'sd5;
        fc1_weights[23][104] = 16'sd31;
        fc1_weights[23][105] = 16'sd-52;
        fc1_weights[23][106] = 16'sd30;
        fc1_weights[23][107] = 16'sd9;
        fc1_weights[23][108] = 16'sd-18;
        fc1_weights[23][109] = 16'sd72;
        fc1_weights[23][110] = 16'sd25;
        fc1_weights[23][111] = 16'sd39;
        fc1_weights[23][112] = 16'sd31;
        fc1_weights[23][113] = 16'sd-54;
        fc1_weights[23][114] = 16'sd14;
        fc1_weights[23][115] = 16'sd-17;
        fc1_weights[23][116] = 16'sd29;
        fc1_weights[23][117] = 16'sd15;
        fc1_weights[23][118] = 16'sd30;
        fc1_weights[23][119] = 16'sd-23;
        fc1_weights[23][120] = 16'sd-38;
        fc1_weights[23][121] = 16'sd8;
        fc1_weights[23][122] = 16'sd-6;
        fc1_weights[23][123] = 16'sd-45;
        fc1_weights[23][124] = 16'sd-4;
        fc1_weights[23][125] = 16'sd-7;
        fc1_weights[23][126] = 16'sd20;
        fc1_weights[23][127] = 16'sd35;
        fc1_weights[23][128] = 16'sd7;
        fc1_weights[23][129] = 16'sd18;
        fc1_weights[23][130] = 16'sd-6;
        fc1_weights[23][131] = 16'sd48;
        fc1_weights[23][132] = 16'sd36;
        fc1_weights[23][133] = 16'sd6;
        fc1_weights[23][134] = 16'sd5;
        fc1_weights[23][135] = 16'sd74;
        fc1_weights[23][136] = 16'sd59;
        fc1_weights[23][137] = 16'sd19;
        fc1_weights[23][138] = 16'sd53;
        fc1_weights[23][139] = 16'sd-49;
        fc1_weights[23][140] = 16'sd-7;
        fc1_weights[23][141] = 16'sd65;
        fc1_weights[23][142] = 16'sd-40;
        fc1_weights[23][143] = 16'sd30;
        fc1_weights[23][144] = 16'sd88;
        fc1_weights[23][145] = 16'sd38;
        fc1_weights[23][146] = 16'sd17;
        fc1_weights[23][147] = 16'sd13;
        fc1_weights[23][148] = 16'sd-44;
        fc1_weights[23][149] = 16'sd-27;
        fc1_weights[23][150] = 16'sd29;
        fc1_weights[23][151] = 16'sd52;
        fc1_weights[23][152] = 16'sd11;
        fc1_weights[23][153] = 16'sd-31;
        fc1_weights[23][154] = 16'sd40;
        fc1_weights[23][155] = 16'sd-39;
        fc1_weights[23][156] = 16'sd-4;
        fc1_weights[23][157] = 16'sd21;
        fc1_weights[23][158] = 16'sd19;
        fc1_weights[23][159] = 16'sd73;
        fc1_weights[23][160] = 16'sd-6;
        fc1_weights[23][161] = 16'sd59;
        fc1_weights[23][162] = 16'sd42;
        fc1_weights[23][163] = 16'sd14;
        fc1_weights[23][164] = 16'sd12;
        fc1_weights[23][165] = 16'sd-5;
        fc1_weights[23][166] = 16'sd-35;
        fc1_weights[23][167] = 16'sd-16;
        fc1_weights[23][168] = 16'sd-25;
        fc1_weights[23][169] = 16'sd38;
        fc1_weights[23][170] = 16'sd25;
        fc1_weights[23][171] = 16'sd-47;
        fc1_weights[23][172] = 16'sd13;
        fc1_weights[23][173] = 16'sd-45;
        fc1_weights[23][174] = 16'sd7;
        fc1_weights[23][175] = 16'sd-35;
        fc1_weights[23][176] = 16'sd-23;
        fc1_weights[23][177] = 16'sd-26;
        fc1_weights[23][178] = 16'sd48;
        fc1_weights[23][179] = 16'sd-2;
        fc1_weights[23][180] = 16'sd28;
        fc1_weights[23][181] = 16'sd52;
        fc1_weights[23][182] = 16'sd58;
        fc1_weights[23][183] = 16'sd41;
        fc1_weights[23][184] = 16'sd66;
        fc1_weights[23][185] = 16'sd-1;
        fc1_weights[23][186] = 16'sd-27;
        fc1_weights[23][187] = 16'sd-50;
        fc1_weights[23][188] = 16'sd-6;
        fc1_weights[23][189] = 16'sd19;
        fc1_weights[23][190] = 16'sd26;
        fc1_weights[23][191] = 16'sd8;
        fc1_weights[23][192] = 16'sd49;
        fc1_weights[23][193] = 16'sd36;
        fc1_weights[23][194] = 16'sd20;
        fc1_weights[23][195] = 16'sd23;
        fc1_weights[23][196] = 16'sd21;
        fc1_weights[23][197] = 16'sd22;
        fc1_weights[23][198] = 16'sd-32;
        fc1_weights[23][199] = 16'sd-32;
        fc1_weights[23][200] = 16'sd43;
        fc1_weights[23][201] = 16'sd-35;
        fc1_weights[23][202] = 16'sd-17;
        fc1_weights[23][203] = 16'sd36;
        fc1_weights[23][204] = 16'sd0;
        fc1_weights[23][205] = 16'sd-23;
        fc1_weights[23][206] = 16'sd13;
        fc1_weights[23][207] = 16'sd62;
        fc1_weights[24][0] = 16'sd-8;
        fc1_weights[24][1] = 16'sd-21;
        fc1_weights[24][2] = 16'sd-29;
        fc1_weights[24][3] = 16'sd16;
        fc1_weights[24][4] = 16'sd-32;
        fc1_weights[24][5] = 16'sd-4;
        fc1_weights[24][6] = 16'sd6;
        fc1_weights[24][7] = 16'sd58;
        fc1_weights[24][8] = 16'sd1;
        fc1_weights[24][9] = 16'sd1;
        fc1_weights[24][10] = 16'sd100;
        fc1_weights[24][11] = 16'sd80;
        fc1_weights[24][12] = 16'sd-24;
        fc1_weights[24][13] = 16'sd-74;
        fc1_weights[24][14] = 16'sd-21;
        fc1_weights[24][15] = 16'sd14;
        fc1_weights[24][16] = 16'sd29;
        fc1_weights[24][17] = 16'sd-6;
        fc1_weights[24][18] = 16'sd-4;
        fc1_weights[24][19] = 16'sd-6;
        fc1_weights[24][20] = 16'sd-4;
        fc1_weights[24][21] = 16'sd-5;
        fc1_weights[24][22] = 16'sd1;
        fc1_weights[24][23] = 16'sd-11;
        fc1_weights[24][24] = 16'sd-2;
        fc1_weights[24][25] = 16'sd-15;
        fc1_weights[24][26] = 16'sd-20;
        fc1_weights[24][27] = 16'sd-28;
        fc1_weights[24][28] = 16'sd2;
        fc1_weights[24][29] = 16'sd44;
        fc1_weights[24][30] = 16'sd14;
        fc1_weights[24][31] = 16'sd25;
        fc1_weights[24][32] = 16'sd-5;
        fc1_weights[24][33] = 16'sd-43;
        fc1_weights[24][34] = 16'sd5;
        fc1_weights[24][35] = 16'sd-33;
        fc1_weights[24][36] = 16'sd43;
        fc1_weights[24][37] = 16'sd123;
        fc1_weights[24][38] = 16'sd25;
        fc1_weights[24][39] = 16'sd-38;
        fc1_weights[24][40] = 16'sd54;
        fc1_weights[24][41] = 16'sd-14;
        fc1_weights[24][42] = 16'sd-12;
        fc1_weights[24][43] = 16'sd86;
        fc1_weights[24][44] = 16'sd53;
        fc1_weights[24][45] = 16'sd-3;
        fc1_weights[24][46] = 16'sd-26;
        fc1_weights[24][47] = 16'sd-58;
        fc1_weights[24][48] = 16'sd14;
        fc1_weights[24][49] = 16'sd-26;
        fc1_weights[24][50] = 16'sd-43;
        fc1_weights[24][51] = 16'sd-50;
        fc1_weights[24][52] = 16'sd-79;
        fc1_weights[24][53] = 16'sd-19;
        fc1_weights[24][54] = 16'sd6;
        fc1_weights[24][55] = 16'sd-21;
        fc1_weights[24][56] = 16'sd-7;
        fc1_weights[24][57] = 16'sd40;
        fc1_weights[24][58] = 16'sd-43;
        fc1_weights[24][59] = 16'sd-57;
        fc1_weights[24][60] = 16'sd-3;
        fc1_weights[24][61] = 16'sd-1;
        fc1_weights[24][62] = 16'sd3;
        fc1_weights[24][63] = 16'sd-16;
        fc1_weights[24][64] = 16'sd-2;
        fc1_weights[24][65] = 16'sd19;
        fc1_weights[24][66] = 16'sd11;
        fc1_weights[24][67] = 16'sd20;
        fc1_weights[24][68] = 16'sd13;
        fc1_weights[24][69] = 16'sd63;
        fc1_weights[24][70] = 16'sd22;
        fc1_weights[24][71] = 16'sd-2;
        fc1_weights[24][72] = 16'sd16;
        fc1_weights[24][73] = 16'sd-8;
        fc1_weights[24][74] = 16'sd9;
        fc1_weights[24][75] = 16'sd-37;
        fc1_weights[24][76] = 16'sd24;
        fc1_weights[24][77] = 16'sd19;
        fc1_weights[24][78] = 16'sd8;
        fc1_weights[24][79] = 16'sd3;
        fc1_weights[24][80] = 16'sd-19;
        fc1_weights[24][81] = 16'sd-14;
        fc1_weights[24][82] = 16'sd-10;
        fc1_weights[24][83] = 16'sd-36;
        fc1_weights[24][84] = 16'sd1;
        fc1_weights[24][85] = 16'sd-46;
        fc1_weights[24][86] = 16'sd-13;
        fc1_weights[24][87] = 16'sd8;
        fc1_weights[24][88] = 16'sd-6;
        fc1_weights[24][89] = 16'sd25;
        fc1_weights[24][90] = 16'sd35;
        fc1_weights[24][91] = 16'sd27;
        fc1_weights[24][92] = 16'sd11;
        fc1_weights[24][93] = 16'sd38;
        fc1_weights[24][94] = 16'sd33;
        fc1_weights[24][95] = 16'sd5;
        fc1_weights[24][96] = 16'sd-14;
        fc1_weights[24][97] = 16'sd23;
        fc1_weights[24][98] = 16'sd-2;
        fc1_weights[24][99] = 16'sd0;
        fc1_weights[24][100] = 16'sd33;
        fc1_weights[24][101] = 16'sd54;
        fc1_weights[24][102] = 16'sd35;
        fc1_weights[24][103] = 16'sd4;
        fc1_weights[24][104] = 16'sd-42;
        fc1_weights[24][105] = 16'sd-29;
        fc1_weights[24][106] = 16'sd-34;
        fc1_weights[24][107] = 16'sd-19;
        fc1_weights[24][108] = 16'sd-21;
        fc1_weights[24][109] = 16'sd-5;
        fc1_weights[24][110] = 16'sd-8;
        fc1_weights[24][111] = 16'sd-29;
        fc1_weights[24][112] = 16'sd20;
        fc1_weights[24][113] = 16'sd8;
        fc1_weights[24][114] = 16'sd-12;
        fc1_weights[24][115] = 16'sd-5;
        fc1_weights[24][116] = 16'sd56;
        fc1_weights[24][117] = 16'sd0;
        fc1_weights[24][118] = 16'sd-46;
        fc1_weights[24][119] = 16'sd22;
        fc1_weights[24][120] = 16'sd-13;
        fc1_weights[24][121] = 16'sd-15;
        fc1_weights[24][122] = 16'sd15;
        fc1_weights[24][123] = 16'sd3;
        fc1_weights[24][124] = 16'sd-5;
        fc1_weights[24][125] = 16'sd-5;
        fc1_weights[24][126] = 16'sd-12;
        fc1_weights[24][127] = 16'sd9;
        fc1_weights[24][128] = 16'sd42;
        fc1_weights[24][129] = 16'sd22;
        fc1_weights[24][130] = 16'sd1;
        fc1_weights[24][131] = 16'sd-24;
        fc1_weights[24][132] = 16'sd3;
        fc1_weights[24][133] = 16'sd-16;
        fc1_weights[24][134] = 16'sd-8;
        fc1_weights[24][135] = 16'sd2;
        fc1_weights[24][136] = 16'sd30;
        fc1_weights[24][137] = 16'sd-15;
        fc1_weights[24][138] = 16'sd100;
        fc1_weights[24][139] = 16'sd45;
        fc1_weights[24][140] = 16'sd-2;
        fc1_weights[24][141] = 16'sd-7;
        fc1_weights[24][142] = 16'sd34;
        fc1_weights[24][143] = 16'sd-11;
        fc1_weights[24][144] = 16'sd40;
        fc1_weights[24][145] = 16'sd19;
        fc1_weights[24][146] = 16'sd35;
        fc1_weights[24][147] = 16'sd-33;
        fc1_weights[24][148] = 16'sd58;
        fc1_weights[24][149] = 16'sd47;
        fc1_weights[24][150] = 16'sd-16;
        fc1_weights[24][151] = 16'sd-23;
        fc1_weights[24][152] = 16'sd7;
        fc1_weights[24][153] = 16'sd-4;
        fc1_weights[24][154] = 16'sd-5;
        fc1_weights[24][155] = 16'sd28;
        fc1_weights[24][156] = 16'sd-14;
        fc1_weights[24][157] = 16'sd-33;
        fc1_weights[24][158] = 16'sd-8;
        fc1_weights[24][159] = 16'sd16;
        fc1_weights[24][160] = 16'sd-6;
        fc1_weights[24][161] = 16'sd-39;
        fc1_weights[24][162] = 16'sd52;
        fc1_weights[24][163] = 16'sd-18;
        fc1_weights[24][164] = 16'sd-9;
        fc1_weights[24][165] = 16'sd16;
        fc1_weights[24][166] = 16'sd29;
        fc1_weights[24][167] = 16'sd24;
        fc1_weights[24][168] = 16'sd50;
        fc1_weights[24][169] = 16'sd-5;
        fc1_weights[24][170] = 16'sd-8;
        fc1_weights[24][171] = 16'sd32;
        fc1_weights[24][172] = 16'sd24;
        fc1_weights[24][173] = 16'sd-6;
        fc1_weights[24][174] = 16'sd16;
        fc1_weights[24][175] = 16'sd-4;
        fc1_weights[24][176] = 16'sd6;
        fc1_weights[24][177] = 16'sd67;
        fc1_weights[24][178] = 16'sd-5;
        fc1_weights[24][179] = 16'sd45;
        fc1_weights[24][180] = 16'sd39;
        fc1_weights[24][181] = 16'sd22;
        fc1_weights[24][182] = 16'sd-2;
        fc1_weights[24][183] = 16'sd7;
        fc1_weights[24][184] = 16'sd-35;
        fc1_weights[24][185] = 16'sd35;
        fc1_weights[24][186] = 16'sd-24;
        fc1_weights[24][187] = 16'sd-20;
        fc1_weights[24][188] = 16'sd7;
        fc1_weights[24][189] = 16'sd-66;
        fc1_weights[24][190] = 16'sd5;
        fc1_weights[24][191] = 16'sd47;
        fc1_weights[24][192] = 16'sd-26;
        fc1_weights[24][193] = 16'sd-7;
        fc1_weights[24][194] = 16'sd0;
        fc1_weights[24][195] = 16'sd-25;
        fc1_weights[24][196] = 16'sd-54;
        fc1_weights[24][197] = 16'sd32;
        fc1_weights[24][198] = 16'sd38;
        fc1_weights[24][199] = 16'sd-19;
        fc1_weights[24][200] = 16'sd5;
        fc1_weights[24][201] = 16'sd-9;
        fc1_weights[24][202] = 16'sd-1;
        fc1_weights[24][203] = 16'sd-13;
        fc1_weights[24][204] = 16'sd50;
        fc1_weights[24][205] = 16'sd30;
        fc1_weights[24][206] = 16'sd10;
        fc1_weights[24][207] = 16'sd11;
        fc1_weights[25][0] = 16'sd-17;
        fc1_weights[25][1] = 16'sd-2;
        fc1_weights[25][2] = 16'sd-1;
        fc1_weights[25][3] = 16'sd30;
        fc1_weights[25][4] = 16'sd-6;
        fc1_weights[25][5] = 16'sd-21;
        fc1_weights[25][6] = 16'sd-2;
        fc1_weights[25][7] = 16'sd27;
        fc1_weights[25][8] = 16'sd12;
        fc1_weights[25][9] = 16'sd-23;
        fc1_weights[25][10] = 16'sd-7;
        fc1_weights[25][11] = 16'sd-1;
        fc1_weights[25][12] = 16'sd-59;
        fc1_weights[25][13] = 16'sd-31;
        fc1_weights[25][14] = 16'sd-4;
        fc1_weights[25][15] = 16'sd2;
        fc1_weights[25][16] = 16'sd-26;
        fc1_weights[25][17] = 16'sd16;
        fc1_weights[25][18] = 16'sd9;
        fc1_weights[25][19] = 16'sd-6;
        fc1_weights[25][20] = 16'sd-4;
        fc1_weights[25][21] = 16'sd-6;
        fc1_weights[25][22] = 16'sd-31;
        fc1_weights[25][23] = 16'sd28;
        fc1_weights[25][24] = 16'sd3;
        fc1_weights[25][25] = 16'sd28;
        fc1_weights[25][26] = 16'sd9;
        fc1_weights[25][27] = 16'sd25;
        fc1_weights[25][28] = 16'sd-9;
        fc1_weights[25][29] = 16'sd42;
        fc1_weights[25][30] = 16'sd41;
        fc1_weights[25][31] = 16'sd20;
        fc1_weights[25][32] = 16'sd23;
        fc1_weights[25][33] = 16'sd-11;
        fc1_weights[25][34] = 16'sd43;
        fc1_weights[25][35] = 16'sd37;
        fc1_weights[25][36] = 16'sd20;
        fc1_weights[25][37] = 16'sd66;
        fc1_weights[25][38] = 16'sd-15;
        fc1_weights[25][39] = 16'sd-27;
        fc1_weights[25][40] = 16'sd-1;
        fc1_weights[25][41] = 16'sd-2;
        fc1_weights[25][42] = 16'sd31;
        fc1_weights[25][43] = 16'sd5;
        fc1_weights[25][44] = 16'sd-4;
        fc1_weights[25][45] = 16'sd-49;
        fc1_weights[25][46] = 16'sd-54;
        fc1_weights[25][47] = 16'sd-74;
        fc1_weights[25][48] = 16'sd-19;
        fc1_weights[25][49] = 16'sd43;
        fc1_weights[25][50] = 16'sd24;
        fc1_weights[25][51] = 16'sd-11;
        fc1_weights[25][52] = 16'sd26;
        fc1_weights[25][53] = 16'sd17;
        fc1_weights[25][54] = 16'sd13;
        fc1_weights[25][55] = 16'sd42;
        fc1_weights[25][56] = 16'sd55;
        fc1_weights[25][57] = 16'sd32;
        fc1_weights[25][58] = 16'sd25;
        fc1_weights[25][59] = 16'sd3;
        fc1_weights[25][60] = 16'sd-26;
        fc1_weights[25][61] = 16'sd0;
        fc1_weights[25][62] = 16'sd10;
        fc1_weights[25][63] = 16'sd25;
        fc1_weights[25][64] = 16'sd1;
        fc1_weights[25][65] = 16'sd-63;
        fc1_weights[25][66] = 16'sd-7;
        fc1_weights[25][67] = 16'sd-45;
        fc1_weights[25][68] = 16'sd-5;
        fc1_weights[25][69] = 16'sd-13;
        fc1_weights[25][70] = 16'sd-3;
        fc1_weights[25][71] = 16'sd-49;
        fc1_weights[25][72] = 16'sd-49;
        fc1_weights[25][73] = 16'sd-41;
        fc1_weights[25][74] = 16'sd-12;
        fc1_weights[25][75] = 16'sd21;
        fc1_weights[25][76] = 16'sd28;
        fc1_weights[25][77] = 16'sd-2;
        fc1_weights[25][78] = 16'sd29;
        fc1_weights[25][79] = 16'sd-10;
        fc1_weights[25][80] = 16'sd-4;
        fc1_weights[25][81] = 16'sd-17;
        fc1_weights[25][82] = 16'sd-3;
        fc1_weights[25][83] = 16'sd-1;
        fc1_weights[25][84] = 16'sd-14;
        fc1_weights[25][85] = 16'sd-62;
        fc1_weights[25][86] = 16'sd-18;
        fc1_weights[25][87] = 16'sd18;
        fc1_weights[25][88] = 16'sd-54;
        fc1_weights[25][89] = 16'sd-39;
        fc1_weights[25][90] = 16'sd-19;
        fc1_weights[25][91] = 16'sd-16;
        fc1_weights[25][92] = 16'sd17;
        fc1_weights[25][93] = 16'sd36;
        fc1_weights[25][94] = 16'sd20;
        fc1_weights[25][95] = 16'sd-1;
        fc1_weights[25][96] = 16'sd-21;
        fc1_weights[25][97] = 16'sd-6;
        fc1_weights[25][98] = 16'sd-18;
        fc1_weights[25][99] = 16'sd4;
        fc1_weights[25][100] = 16'sd-3;
        fc1_weights[25][101] = 16'sd37;
        fc1_weights[25][102] = 16'sd35;
        fc1_weights[25][103] = 16'sd36;
        fc1_weights[25][104] = 16'sd3;
        fc1_weights[25][105] = 16'sd-13;
        fc1_weights[25][106] = 16'sd8;
        fc1_weights[25][107] = 16'sd-31;
        fc1_weights[25][108] = 16'sd3;
        fc1_weights[25][109] = 16'sd-8;
        fc1_weights[25][110] = 16'sd-35;
        fc1_weights[25][111] = 16'sd-11;
        fc1_weights[25][112] = 16'sd-13;
        fc1_weights[25][113] = 16'sd7;
        fc1_weights[25][114] = 16'sd-37;
        fc1_weights[25][115] = 16'sd-10;
        fc1_weights[25][116] = 16'sd-58;
        fc1_weights[25][117] = 16'sd8;
        fc1_weights[25][118] = 16'sd21;
        fc1_weights[25][119] = 16'sd22;
        fc1_weights[25][120] = 16'sd-36;
        fc1_weights[25][121] = 16'sd-17;
        fc1_weights[25][122] = 16'sd-43;
        fc1_weights[25][123] = 16'sd12;
        fc1_weights[25][124] = 16'sd-1;
        fc1_weights[25][125] = 16'sd-46;
        fc1_weights[25][126] = 16'sd-37;
        fc1_weights[25][127] = 16'sd-5;
        fc1_weights[25][128] = 16'sd35;
        fc1_weights[25][129] = 16'sd-9;
        fc1_weights[25][130] = 16'sd-24;
        fc1_weights[25][131] = 16'sd-44;
        fc1_weights[25][132] = 16'sd-41;
        fc1_weights[25][133] = 16'sd-31;
        fc1_weights[25][134] = 16'sd-7;
        fc1_weights[25][135] = 16'sd-6;
        fc1_weights[25][136] = 16'sd-21;
        fc1_weights[25][137] = 16'sd5;
        fc1_weights[25][138] = 16'sd37;
        fc1_weights[25][139] = 16'sd45;
        fc1_weights[25][140] = 16'sd61;
        fc1_weights[25][141] = 16'sd32;
        fc1_weights[25][142] = 16'sd51;
        fc1_weights[25][143] = 16'sd62;
        fc1_weights[25][144] = 16'sd42;
        fc1_weights[25][145] = 16'sd23;
        fc1_weights[25][146] = 16'sd20;
        fc1_weights[25][147] = 16'sd47;
        fc1_weights[25][148] = 16'sd59;
        fc1_weights[25][149] = 16'sd36;
        fc1_weights[25][150] = 16'sd30;
        fc1_weights[25][151] = 16'sd9;
        fc1_weights[25][152] = 16'sd-4;
        fc1_weights[25][153] = 16'sd1;
        fc1_weights[25][154] = 16'sd0;
        fc1_weights[25][155] = 16'sd-14;
        fc1_weights[25][156] = 16'sd14;
        fc1_weights[25][157] = 16'sd4;
        fc1_weights[25][158] = 16'sd-39;
        fc1_weights[25][159] = 16'sd-75;
        fc1_weights[25][160] = 16'sd26;
        fc1_weights[25][161] = 16'sd-6;
        fc1_weights[25][162] = 16'sd58;
        fc1_weights[25][163] = 16'sd42;
        fc1_weights[25][164] = 16'sd42;
        fc1_weights[25][165] = 16'sd46;
        fc1_weights[25][166] = 16'sd18;
        fc1_weights[25][167] = 16'sd6;
        fc1_weights[25][168] = 16'sd48;
        fc1_weights[25][169] = 16'sd33;
        fc1_weights[25][170] = 16'sd19;
        fc1_weights[25][171] = 16'sd9;
        fc1_weights[25][172] = 16'sd31;
        fc1_weights[25][173] = 16'sd-5;
        fc1_weights[25][174] = 16'sd-7;
        fc1_weights[25][175] = 16'sd-13;
        fc1_weights[25][176] = 16'sd8;
        fc1_weights[25][177] = 16'sd2;
        fc1_weights[25][178] = 16'sd-31;
        fc1_weights[25][179] = 16'sd15;
        fc1_weights[25][180] = 16'sd-4;
        fc1_weights[25][181] = 16'sd-1;
        fc1_weights[25][182] = 16'sd12;
        fc1_weights[25][183] = 16'sd-12;
        fc1_weights[25][184] = 16'sd-23;
        fc1_weights[25][185] = 16'sd-1;
        fc1_weights[25][186] = 16'sd72;
        fc1_weights[25][187] = 16'sd28;
        fc1_weights[25][188] = 16'sd35;
        fc1_weights[25][189] = 16'sd36;
        fc1_weights[25][190] = 16'sd27;
        fc1_weights[25][191] = 16'sd-14;
        fc1_weights[25][192] = 16'sd-5;
        fc1_weights[25][193] = 16'sd-13;
        fc1_weights[25][194] = 16'sd1;
        fc1_weights[25][195] = 16'sd17;
        fc1_weights[25][196] = 16'sd18;
        fc1_weights[25][197] = 16'sd8;
        fc1_weights[25][198] = 16'sd-18;
        fc1_weights[25][199] = 16'sd17;
        fc1_weights[25][200] = 16'sd11;
        fc1_weights[25][201] = 16'sd3;
        fc1_weights[25][202] = 16'sd-17;
        fc1_weights[25][203] = 16'sd41;
        fc1_weights[25][204] = 16'sd34;
        fc1_weights[25][205] = 16'sd4;
        fc1_weights[25][206] = 16'sd-1;
        fc1_weights[25][207] = 16'sd-4;
        fc1_weights[26][0] = 16'sd19;
        fc1_weights[26][1] = 16'sd-9;
        fc1_weights[26][2] = 16'sd-7;
        fc1_weights[26][3] = 16'sd47;
        fc1_weights[26][4] = 16'sd25;
        fc1_weights[26][5] = 16'sd46;
        fc1_weights[26][6] = 16'sd28;
        fc1_weights[26][7] = 16'sd-43;
        fc1_weights[26][8] = 16'sd16;
        fc1_weights[26][9] = 16'sd-13;
        fc1_weights[26][10] = 16'sd-4;
        fc1_weights[26][11] = 16'sd13;
        fc1_weights[26][12] = 16'sd-29;
        fc1_weights[26][13] = 16'sd-47;
        fc1_weights[26][14] = 16'sd-12;
        fc1_weights[26][15] = 16'sd22;
        fc1_weights[26][16] = 16'sd6;
        fc1_weights[26][17] = 16'sd-24;
        fc1_weights[26][18] = 16'sd-41;
        fc1_weights[26][19] = 16'sd5;
        fc1_weights[26][20] = 16'sd-10;
        fc1_weights[26][21] = 16'sd-31;
        fc1_weights[26][22] = 16'sd-18;
        fc1_weights[26][23] = 16'sd-52;
        fc1_weights[26][24] = 16'sd-7;
        fc1_weights[26][25] = 16'sd-23;
        fc1_weights[26][26] = 16'sd-4;
        fc1_weights[26][27] = 16'sd23;
        fc1_weights[26][28] = 16'sd2;
        fc1_weights[26][29] = 16'sd4;
        fc1_weights[26][30] = 16'sd25;
        fc1_weights[26][31] = 16'sd18;
        fc1_weights[26][32] = 16'sd33;
        fc1_weights[26][33] = 16'sd-9;
        fc1_weights[26][34] = 16'sd-11;
        fc1_weights[26][35] = 16'sd-11;
        fc1_weights[26][36] = 16'sd25;
        fc1_weights[26][37] = 16'sd-54;
        fc1_weights[26][38] = 16'sd-37;
        fc1_weights[26][39] = 16'sd9;
        fc1_weights[26][40] = 16'sd20;
        fc1_weights[26][41] = 16'sd33;
        fc1_weights[26][42] = 16'sd-8;
        fc1_weights[26][43] = 16'sd57;
        fc1_weights[26][44] = 16'sd38;
        fc1_weights[26][45] = 16'sd52;
        fc1_weights[26][46] = 16'sd43;
        fc1_weights[26][47] = 16'sd-2;
        fc1_weights[26][48] = 16'sd-17;
        fc1_weights[26][49] = 16'sd-1;
        fc1_weights[26][50] = 16'sd-17;
        fc1_weights[26][51] = 16'sd14;
        fc1_weights[26][52] = 16'sd-19;
        fc1_weights[26][53] = 16'sd30;
        fc1_weights[26][54] = 16'sd30;
        fc1_weights[26][55] = 16'sd25;
        fc1_weights[26][56] = 16'sd22;
        fc1_weights[26][57] = 16'sd18;
        fc1_weights[26][58] = 16'sd-10;
        fc1_weights[26][59] = 16'sd-10;
        fc1_weights[26][60] = 16'sd2;
        fc1_weights[26][61] = 16'sd-14;
        fc1_weights[26][62] = 16'sd32;
        fc1_weights[26][63] = 16'sd0;
        fc1_weights[26][64] = 16'sd-11;
        fc1_weights[26][65] = 16'sd-1;
        fc1_weights[26][66] = 16'sd4;
        fc1_weights[26][67] = 16'sd-11;
        fc1_weights[26][68] = 16'sd-34;
        fc1_weights[26][69] = 16'sd17;
        fc1_weights[26][70] = 16'sd6;
        fc1_weights[26][71] = 16'sd-10;
        fc1_weights[26][72] = 16'sd-33;
        fc1_weights[26][73] = 16'sd-43;
        fc1_weights[26][74] = 16'sd-21;
        fc1_weights[26][75] = 16'sd-35;
        fc1_weights[26][76] = 16'sd-17;
        fc1_weights[26][77] = 16'sd-9;
        fc1_weights[26][78] = 16'sd3;
        fc1_weights[26][79] = 16'sd10;
        fc1_weights[26][80] = 16'sd-6;
        fc1_weights[26][81] = 16'sd1;
        fc1_weights[26][82] = 16'sd29;
        fc1_weights[26][83] = 16'sd1;
        fc1_weights[26][84] = 16'sd-40;
        fc1_weights[26][85] = 16'sd-9;
        fc1_weights[26][86] = 16'sd-7;
        fc1_weights[26][87] = 16'sd13;
        fc1_weights[26][88] = 16'sd21;
        fc1_weights[26][89] = 16'sd5;
        fc1_weights[26][90] = 16'sd-1;
        fc1_weights[26][91] = 16'sd-11;
        fc1_weights[26][92] = 16'sd-17;
        fc1_weights[26][93] = 16'sd-5;
        fc1_weights[26][94] = 16'sd3;
        fc1_weights[26][95] = 16'sd22;
        fc1_weights[26][96] = 16'sd5;
        fc1_weights[26][97] = 16'sd10;
        fc1_weights[26][98] = 16'sd-32;
        fc1_weights[26][99] = 16'sd-14;
        fc1_weights[26][100] = 16'sd-21;
        fc1_weights[26][101] = 16'sd-16;
        fc1_weights[26][102] = 16'sd-9;
        fc1_weights[26][103] = 16'sd-27;
        fc1_weights[26][104] = 16'sd3;
        fc1_weights[26][105] = 16'sd28;
        fc1_weights[26][106] = 16'sd15;
        fc1_weights[26][107] = 16'sd27;
        fc1_weights[26][108] = 16'sd18;
        fc1_weights[26][109] = 16'sd10;
        fc1_weights[26][110] = 16'sd-8;
        fc1_weights[26][111] = 16'sd7;
        fc1_weights[26][112] = 16'sd22;
        fc1_weights[26][113] = 16'sd-3;
        fc1_weights[26][114] = 16'sd-4;
        fc1_weights[26][115] = 16'sd7;
        fc1_weights[26][116] = 16'sd17;
        fc1_weights[26][117] = 16'sd11;
        fc1_weights[26][118] = 16'sd-27;
        fc1_weights[26][119] = 16'sd11;
        fc1_weights[26][120] = 16'sd12;
        fc1_weights[26][121] = 16'sd4;
        fc1_weights[26][122] = 16'sd7;
        fc1_weights[26][123] = 16'sd30;
        fc1_weights[26][124] = 16'sd-27;
        fc1_weights[26][125] = 16'sd-15;
        fc1_weights[26][126] = 16'sd8;
        fc1_weights[26][127] = 16'sd-20;
        fc1_weights[26][128] = 16'sd-11;
        fc1_weights[26][129] = 16'sd-25;
        fc1_weights[26][130] = 16'sd-4;
        fc1_weights[26][131] = 16'sd12;
        fc1_weights[26][132] = 16'sd1;
        fc1_weights[26][133] = 16'sd-10;
        fc1_weights[26][134] = 16'sd17;
        fc1_weights[26][135] = 16'sd28;
        fc1_weights[26][136] = 16'sd-8;
        fc1_weights[26][137] = 16'sd32;
        fc1_weights[26][138] = 16'sd-31;
        fc1_weights[26][139] = 16'sd-9;
        fc1_weights[26][140] = 16'sd-32;
        fc1_weights[26][141] = 16'sd-52;
        fc1_weights[26][142] = 16'sd-17;
        fc1_weights[26][143] = 16'sd-35;
        fc1_weights[26][144] = 16'sd-8;
        fc1_weights[26][145] = 16'sd-55;
        fc1_weights[26][146] = 16'sd-16;
        fc1_weights[26][147] = 16'sd-25;
        fc1_weights[26][148] = 16'sd-33;
        fc1_weights[26][149] = 16'sd-11;
        fc1_weights[26][150] = 16'sd-29;
        fc1_weights[26][151] = 16'sd-9;
        fc1_weights[26][152] = 16'sd-22;
        fc1_weights[26][153] = 16'sd-10;
        fc1_weights[26][154] = 16'sd-3;
        fc1_weights[26][155] = 16'sd-8;
        fc1_weights[26][156] = 16'sd-3;
        fc1_weights[26][157] = 16'sd-6;
        fc1_weights[26][158] = 16'sd2;
        fc1_weights[26][159] = 16'sd0;
        fc1_weights[26][160] = 16'sd-10;
        fc1_weights[26][161] = 16'sd-13;
        fc1_weights[26][162] = 16'sd3;
        fc1_weights[26][163] = 16'sd0;
        fc1_weights[26][164] = 16'sd7;
        fc1_weights[26][165] = 16'sd-15;
        fc1_weights[26][166] = 16'sd-12;
        fc1_weights[26][167] = 16'sd4;
        fc1_weights[26][168] = 16'sd14;
        fc1_weights[26][169] = 16'sd0;
        fc1_weights[26][170] = 16'sd10;
        fc1_weights[26][171] = 16'sd19;
        fc1_weights[26][172] = 16'sd-6;
        fc1_weights[26][173] = 16'sd-27;
        fc1_weights[26][174] = 16'sd-65;
        fc1_weights[26][175] = 16'sd-33;
        fc1_weights[26][176] = 16'sd-19;
        fc1_weights[26][177] = 16'sd1;
        fc1_weights[26][178] = 16'sd-33;
        fc1_weights[26][179] = 16'sd-7;
        fc1_weights[26][180] = 16'sd-33;
        fc1_weights[26][181] = 16'sd-32;
        fc1_weights[26][182] = 16'sd4;
        fc1_weights[26][183] = 16'sd31;
        fc1_weights[26][184] = 16'sd19;
        fc1_weights[26][185] = 16'sd48;
        fc1_weights[26][186] = 16'sd27;
        fc1_weights[26][187] = 16'sd34;
        fc1_weights[26][188] = 16'sd39;
        fc1_weights[26][189] = 16'sd34;
        fc1_weights[26][190] = 16'sd8;
        fc1_weights[26][191] = 16'sd-6;
        fc1_weights[26][192] = 16'sd5;
        fc1_weights[26][193] = 16'sd2;
        fc1_weights[26][194] = 16'sd14;
        fc1_weights[26][195] = 16'sd15;
        fc1_weights[26][196] = 16'sd28;
        fc1_weights[26][197] = 16'sd53;
        fc1_weights[26][198] = 16'sd24;
        fc1_weights[26][199] = 16'sd-12;
        fc1_weights[26][200] = 16'sd2;
        fc1_weights[26][201] = 16'sd-7;
        fc1_weights[26][202] = 16'sd-9;
        fc1_weights[26][203] = 16'sd5;
        fc1_weights[26][204] = 16'sd-21;
        fc1_weights[26][205] = 16'sd8;
        fc1_weights[26][206] = 16'sd-1;
        fc1_weights[26][207] = 16'sd-18;
        fc1_weights[27][0] = 16'sd33;
        fc1_weights[27][1] = 16'sd14;
        fc1_weights[27][2] = 16'sd4;
        fc1_weights[27][3] = 16'sd-27;
        fc1_weights[27][4] = 16'sd6;
        fc1_weights[27][5] = 16'sd-21;
        fc1_weights[27][6] = 16'sd-2;
        fc1_weights[27][7] = 16'sd4;
        fc1_weights[27][8] = 16'sd-4;
        fc1_weights[27][9] = 16'sd39;
        fc1_weights[27][10] = 16'sd5;
        fc1_weights[27][11] = 16'sd5;
        fc1_weights[27][12] = 16'sd-19;
        fc1_weights[27][13] = 16'sd-27;
        fc1_weights[27][14] = 16'sd-16;
        fc1_weights[27][15] = 16'sd-27;
        fc1_weights[27][16] = 16'sd-31;
        fc1_weights[27][17] = 16'sd-12;
        fc1_weights[27][18] = 16'sd11;
        fc1_weights[27][19] = 16'sd16;
        fc1_weights[27][20] = 16'sd39;
        fc1_weights[27][21] = 16'sd17;
        fc1_weights[27][22] = 16'sd42;
        fc1_weights[27][23] = 16'sd31;
        fc1_weights[27][24] = 16'sd55;
        fc1_weights[27][25] = 16'sd50;
        fc1_weights[27][26] = 16'sd20;
        fc1_weights[27][27] = 16'sd20;
        fc1_weights[27][28] = 16'sd4;
        fc1_weights[27][29] = 16'sd-24;
        fc1_weights[27][30] = 16'sd0;
        fc1_weights[27][31] = 16'sd-29;
        fc1_weights[27][32] = 16'sd-15;
        fc1_weights[27][33] = 16'sd-12;
        fc1_weights[27][34] = 16'sd-2;
        fc1_weights[27][35] = 16'sd23;
        fc1_weights[27][36] = 16'sd44;
        fc1_weights[27][37] = 16'sd-25;
        fc1_weights[27][38] = 16'sd33;
        fc1_weights[27][39] = 16'sd16;
        fc1_weights[27][40] = 16'sd26;
        fc1_weights[27][41] = 16'sd-30;
        fc1_weights[27][42] = 16'sd-16;
        fc1_weights[27][43] = 16'sd19;
        fc1_weights[27][44] = 16'sd-5;
        fc1_weights[27][45] = 16'sd-18;
        fc1_weights[27][46] = 16'sd-8;
        fc1_weights[27][47] = 16'sd42;
        fc1_weights[27][48] = 16'sd40;
        fc1_weights[27][49] = 16'sd18;
        fc1_weights[27][50] = 16'sd42;
        fc1_weights[27][51] = 16'sd17;
        fc1_weights[27][52] = 16'sd30;
        fc1_weights[27][53] = 16'sd21;
        fc1_weights[27][54] = 16'sd16;
        fc1_weights[27][55] = 16'sd23;
        fc1_weights[27][56] = 16'sd2;
        fc1_weights[27][57] = 16'sd2;
        fc1_weights[27][58] = 16'sd-12;
        fc1_weights[27][59] = 16'sd-14;
        fc1_weights[27][60] = 16'sd18;
        fc1_weights[27][61] = 16'sd56;
        fc1_weights[27][62] = 16'sd10;
        fc1_weights[27][63] = 16'sd2;
        fc1_weights[27][64] = 16'sd12;
        fc1_weights[27][65] = 16'sd-20;
        fc1_weights[27][66] = 16'sd-12;
        fc1_weights[27][67] = 16'sd-24;
        fc1_weights[27][68] = 16'sd-20;
        fc1_weights[27][69] = 16'sd-14;
        fc1_weights[27][70] = 16'sd-31;
        fc1_weights[27][71] = 16'sd11;
        fc1_weights[27][72] = 16'sd11;
        fc1_weights[27][73] = 16'sd-4;
        fc1_weights[27][74] = 16'sd6;
        fc1_weights[27][75] = 16'sd18;
        fc1_weights[27][76] = 16'sd32;
        fc1_weights[27][77] = 16'sd10;
        fc1_weights[27][78] = 16'sd25;
        fc1_weights[27][79] = 16'sd57;
        fc1_weights[27][80] = 16'sd-8;
        fc1_weights[27][81] = 16'sd-35;
        fc1_weights[27][82] = 16'sd-33;
        fc1_weights[27][83] = 16'sd-41;
        fc1_weights[27][84] = 16'sd-9;
        fc1_weights[27][85] = 16'sd-23;
        fc1_weights[27][86] = 16'sd3;
        fc1_weights[27][87] = 16'sd36;
        fc1_weights[27][88] = 16'sd2;
        fc1_weights[27][89] = 16'sd2;
        fc1_weights[27][90] = 16'sd16;
        fc1_weights[27][91] = 16'sd-16;
        fc1_weights[27][92] = 16'sd-7;
        fc1_weights[27][93] = 16'sd-29;
        fc1_weights[27][94] = 16'sd-20;
        fc1_weights[27][95] = 16'sd-28;
        fc1_weights[27][96] = 16'sd-43;
        fc1_weights[27][97] = 16'sd-28;
        fc1_weights[27][98] = 16'sd-17;
        fc1_weights[27][99] = 16'sd-20;
        fc1_weights[27][100] = 16'sd22;
        fc1_weights[27][101] = 16'sd31;
        fc1_weights[27][102] = 16'sd-13;
        fc1_weights[27][103] = 16'sd-27;
        fc1_weights[27][104] = 16'sd26;
        fc1_weights[27][105] = 16'sd-18;
        fc1_weights[27][106] = 16'sd-20;
        fc1_weights[27][107] = 16'sd-22;
        fc1_weights[27][108] = 16'sd-2;
        fc1_weights[27][109] = 16'sd-17;
        fc1_weights[27][110] = 16'sd5;
        fc1_weights[27][111] = 16'sd16;
        fc1_weights[27][112] = 16'sd15;
        fc1_weights[27][113] = 16'sd12;
        fc1_weights[27][114] = 16'sd-25;
        fc1_weights[27][115] = 16'sd-16;
        fc1_weights[27][116] = 16'sd-3;
        fc1_weights[27][117] = 16'sd-4;
        fc1_weights[27][118] = 16'sd-26;
        fc1_weights[27][119] = 16'sd-26;
        fc1_weights[27][120] = 16'sd-19;
        fc1_weights[27][121] = 16'sd2;
        fc1_weights[27][122] = 16'sd-29;
        fc1_weights[27][123] = 16'sd7;
        fc1_weights[27][124] = 16'sd-26;
        fc1_weights[27][125] = 16'sd-7;
        fc1_weights[27][126] = 16'sd-60;
        fc1_weights[27][127] = 16'sd4;
        fc1_weights[27][128] = 16'sd-21;
        fc1_weights[27][129] = 16'sd-82;
        fc1_weights[27][130] = 16'sd-2;
        fc1_weights[27][131] = 16'sd7;
        fc1_weights[27][132] = 16'sd-40;
        fc1_weights[27][133] = 16'sd-55;
        fc1_weights[27][134] = 16'sd-25;
        fc1_weights[27][135] = 16'sd-26;
        fc1_weights[27][136] = 16'sd28;
        fc1_weights[27][137] = 16'sd31;
        fc1_weights[27][138] = 16'sd10;
        fc1_weights[27][139] = 16'sd10;
        fc1_weights[27][140] = 16'sd-45;
        fc1_weights[27][141] = 16'sd-32;
        fc1_weights[27][142] = 16'sd-25;
        fc1_weights[27][143] = 16'sd-60;
        fc1_weights[27][144] = 16'sd-30;
        fc1_weights[27][145] = 16'sd-25;
        fc1_weights[27][146] = 16'sd11;
        fc1_weights[27][147] = 16'sd36;
        fc1_weights[27][148] = 16'sd14;
        fc1_weights[27][149] = 16'sd-7;
        fc1_weights[27][150] = 16'sd-15;
        fc1_weights[27][151] = 16'sd-11;
        fc1_weights[27][152] = 16'sd-5;
        fc1_weights[27][153] = 16'sd16;
        fc1_weights[27][154] = 16'sd-36;
        fc1_weights[27][155] = 16'sd-39;
        fc1_weights[27][156] = 16'sd16;
        fc1_weights[27][157] = 16'sd6;
        fc1_weights[27][158] = 16'sd13;
        fc1_weights[27][159] = 16'sd-22;
        fc1_weights[27][160] = 16'sd23;
        fc1_weights[27][161] = 16'sd66;
        fc1_weights[27][162] = 16'sd36;
        fc1_weights[27][163] = 16'sd16;
        fc1_weights[27][164] = 16'sd25;
        fc1_weights[27][165] = 16'sd-30;
        fc1_weights[27][166] = 16'sd-7;
        fc1_weights[27][167] = 16'sd-6;
        fc1_weights[27][168] = 16'sd1;
        fc1_weights[27][169] = 16'sd-1;
        fc1_weights[27][170] = 16'sd3;
        fc1_weights[27][171] = 16'sd-13;
        fc1_weights[27][172] = 16'sd-7;
        fc1_weights[27][173] = 16'sd9;
        fc1_weights[27][174] = 16'sd-3;
        fc1_weights[27][175] = 16'sd-6;
        fc1_weights[27][176] = 16'sd-8;
        fc1_weights[27][177] = 16'sd-11;
        fc1_weights[27][178] = 16'sd-18;
        fc1_weights[27][179] = 16'sd-6;
        fc1_weights[27][180] = 16'sd-30;
        fc1_weights[27][181] = 16'sd-14;
        fc1_weights[27][182] = 16'sd17;
        fc1_weights[27][183] = 16'sd11;
        fc1_weights[27][184] = 16'sd5;
        fc1_weights[27][185] = 16'sd12;
        fc1_weights[27][186] = 16'sd13;
        fc1_weights[27][187] = 16'sd25;
        fc1_weights[27][188] = 16'sd9;
        fc1_weights[27][189] = 16'sd31;
        fc1_weights[27][190] = 16'sd-11;
        fc1_weights[27][191] = 16'sd-11;
        fc1_weights[27][192] = 16'sd-39;
        fc1_weights[27][193] = 16'sd-12;
        fc1_weights[27][194] = 16'sd-2;
        fc1_weights[27][195] = 16'sd-11;
        fc1_weights[27][196] = 16'sd24;
        fc1_weights[27][197] = 16'sd-4;
        fc1_weights[27][198] = 16'sd-19;
        fc1_weights[27][199] = 16'sd-5;
        fc1_weights[27][200] = 16'sd11;
        fc1_weights[27][201] = 16'sd19;
        fc1_weights[27][202] = 16'sd-19;
        fc1_weights[27][203] = 16'sd-5;
        fc1_weights[27][204] = 16'sd-1;
        fc1_weights[27][205] = 16'sd-16;
        fc1_weights[27][206] = 16'sd-11;
        fc1_weights[27][207] = 16'sd-18;
        fc1_weights[28][0] = 16'sd-25;
        fc1_weights[28][1] = 16'sd-65;
        fc1_weights[28][2] = 16'sd-76;
        fc1_weights[28][3] = 16'sd39;
        fc1_weights[28][4] = 16'sd25;
        fc1_weights[28][5] = 16'sd-16;
        fc1_weights[28][6] = 16'sd1;
        fc1_weights[28][7] = 16'sd-36;
        fc1_weights[28][8] = 16'sd66;
        fc1_weights[28][9] = 16'sd26;
        fc1_weights[28][10] = 16'sd-41;
        fc1_weights[28][11] = 16'sd-10;
        fc1_weights[28][12] = 16'sd24;
        fc1_weights[28][13] = 16'sd-27;
        fc1_weights[28][14] = 16'sd-18;
        fc1_weights[28][15] = 16'sd-3;
        fc1_weights[28][16] = 16'sd34;
        fc1_weights[28][17] = 16'sd18;
        fc1_weights[28][18] = 16'sd18;
        fc1_weights[28][19] = 16'sd26;
        fc1_weights[28][20] = 16'sd-11;
        fc1_weights[28][21] = 16'sd-9;
        fc1_weights[28][22] = 16'sd12;
        fc1_weights[28][23] = 16'sd22;
        fc1_weights[28][24] = 16'sd19;
        fc1_weights[28][25] = 16'sd-28;
        fc1_weights[28][26] = 16'sd26;
        fc1_weights[28][27] = 16'sd-54;
        fc1_weights[28][28] = 16'sd-7;
        fc1_weights[28][29] = 16'sd-16;
        fc1_weights[28][30] = 16'sd-28;
        fc1_weights[28][31] = 16'sd-67;
        fc1_weights[28][32] = 16'sd9;
        fc1_weights[28][33] = 16'sd23;
        fc1_weights[28][34] = 16'sd28;
        fc1_weights[28][35] = 16'sd21;
        fc1_weights[28][36] = 16'sd-38;
        fc1_weights[28][37] = 16'sd-80;
        fc1_weights[28][38] = 16'sd-47;
        fc1_weights[28][39] = 16'sd-52;
        fc1_weights[28][40] = 16'sd-45;
        fc1_weights[28][41] = 16'sd-51;
        fc1_weights[28][42] = 16'sd4;
        fc1_weights[28][43] = 16'sd30;
        fc1_weights[28][44] = 16'sd14;
        fc1_weights[28][45] = 16'sd44;
        fc1_weights[28][46] = 16'sd43;
        fc1_weights[28][47] = 16'sd15;
        fc1_weights[28][48] = 16'sd-35;
        fc1_weights[28][49] = 16'sd-1;
        fc1_weights[28][50] = 16'sd-19;
        fc1_weights[28][51] = 16'sd52;
        fc1_weights[28][52] = 16'sd12;
        fc1_weights[28][53] = 16'sd-55;
        fc1_weights[28][54] = 16'sd13;
        fc1_weights[28][55] = 16'sd1;
        fc1_weights[28][56] = 16'sd-3;
        fc1_weights[28][57] = 16'sd-34;
        fc1_weights[28][58] = 16'sd4;
        fc1_weights[28][59] = 16'sd-35;
        fc1_weights[28][60] = 16'sd-44;
        fc1_weights[28][61] = 16'sd-33;
        fc1_weights[28][62] = 16'sd-21;
        fc1_weights[28][63] = 16'sd-88;
        fc1_weights[28][64] = 16'sd-108;
        fc1_weights[28][65] = 16'sd-16;
        fc1_weights[28][66] = 16'sd-31;
        fc1_weights[28][67] = 16'sd-11;
        fc1_weights[28][68] = 16'sd16;
        fc1_weights[28][69] = 16'sd79;
        fc1_weights[28][70] = 16'sd23;
        fc1_weights[28][71] = 16'sd17;
        fc1_weights[28][72] = 16'sd-4;
        fc1_weights[28][73] = 16'sd5;
        fc1_weights[28][74] = 16'sd-26;
        fc1_weights[28][75] = 16'sd-18;
        fc1_weights[28][76] = 16'sd1;
        fc1_weights[28][77] = 16'sd6;
        fc1_weights[28][78] = 16'sd-13;
        fc1_weights[28][79] = 16'sd-19;
        fc1_weights[28][80] = 16'sd2;
        fc1_weights[28][81] = 16'sd38;
        fc1_weights[28][82] = 16'sd39;
        fc1_weights[28][83] = 16'sd20;
        fc1_weights[28][84] = 16'sd29;
        fc1_weights[28][85] = 16'sd17;
        fc1_weights[28][86] = 16'sd11;
        fc1_weights[28][87] = 16'sd39;
        fc1_weights[28][88] = 16'sd33;
        fc1_weights[28][89] = 16'sd-29;
        fc1_weights[28][90] = 16'sd-13;
        fc1_weights[28][91] = 16'sd-18;
        fc1_weights[28][92] = 16'sd-16;
        fc1_weights[28][93] = 16'sd-45;
        fc1_weights[28][94] = 16'sd-13;
        fc1_weights[28][95] = 16'sd-35;
        fc1_weights[28][96] = 16'sd-2;
        fc1_weights[28][97] = 16'sd-13;
        fc1_weights[28][98] = 16'sd-12;
        fc1_weights[28][99] = 16'sd6;
        fc1_weights[28][100] = 16'sd-44;
        fc1_weights[28][101] = 16'sd7;
        fc1_weights[28][102] = 16'sd9;
        fc1_weights[28][103] = 16'sd9;
        fc1_weights[28][104] = 16'sd-15;
        fc1_weights[28][105] = 16'sd0;
        fc1_weights[28][106] = 16'sd12;
        fc1_weights[28][107] = 16'sd49;
        fc1_weights[28][108] = 16'sd-38;
        fc1_weights[28][109] = 16'sd23;
        fc1_weights[28][110] = 16'sd-37;
        fc1_weights[28][111] = 16'sd-43;
        fc1_weights[28][112] = 16'sd22;
        fc1_weights[28][113] = 16'sd58;
        fc1_weights[28][114] = 16'sd8;
        fc1_weights[28][115] = 16'sd22;
        fc1_weights[28][116] = 16'sd31;
        fc1_weights[28][117] = 16'sd26;
        fc1_weights[28][118] = 16'sd-27;
        fc1_weights[28][119] = 16'sd-16;
        fc1_weights[28][120] = 16'sd34;
        fc1_weights[28][121] = 16'sd-11;
        fc1_weights[28][122] = 16'sd-34;
        fc1_weights[28][123] = 16'sd41;
        fc1_weights[28][124] = 16'sd14;
        fc1_weights[28][125] = 16'sd16;
        fc1_weights[28][126] = 16'sd62;
        fc1_weights[28][127] = 16'sd41;
        fc1_weights[28][128] = 16'sd9;
        fc1_weights[28][129] = 16'sd43;
        fc1_weights[28][130] = 16'sd8;
        fc1_weights[28][131] = 16'sd8;
        fc1_weights[28][132] = 16'sd5;
        fc1_weights[28][133] = 16'sd-15;
        fc1_weights[28][134] = 16'sd-45;
        fc1_weights[28][135] = 16'sd-29;
        fc1_weights[28][136] = 16'sd-51;
        fc1_weights[28][137] = 16'sd-56;
        fc1_weights[28][138] = 16'sd-70;
        fc1_weights[28][139] = 16'sd-2;
        fc1_weights[28][140] = 16'sd-27;
        fc1_weights[28][141] = 16'sd-80;
        fc1_weights[28][142] = 16'sd-73;
        fc1_weights[28][143] = 16'sd-36;
        fc1_weights[28][144] = 16'sd8;
        fc1_weights[28][145] = 16'sd49;
        fc1_weights[28][146] = 16'sd28;
        fc1_weights[28][147] = 16'sd-14;
        fc1_weights[28][148] = 16'sd-10;
        fc1_weights[28][149] = 16'sd17;
        fc1_weights[28][150] = 16'sd14;
        fc1_weights[28][151] = 16'sd17;
        fc1_weights[28][152] = 16'sd-24;
        fc1_weights[28][153] = 16'sd-3;
        fc1_weights[28][154] = 16'sd-12;
        fc1_weights[28][155] = 16'sd-19;
        fc1_weights[28][156] = 16'sd21;
        fc1_weights[28][157] = 16'sd-39;
        fc1_weights[28][158] = 16'sd3;
        fc1_weights[28][159] = 16'sd-7;
        fc1_weights[28][160] = 16'sd-13;
        fc1_weights[28][161] = 16'sd5;
        fc1_weights[28][162] = 16'sd-24;
        fc1_weights[28][163] = 16'sd50;
        fc1_weights[28][164] = 16'sd43;
        fc1_weights[28][165] = 16'sd40;
        fc1_weights[28][166] = 16'sd-6;
        fc1_weights[28][167] = 16'sd-5;
        fc1_weights[28][168] = 16'sd-35;
        fc1_weights[28][169] = 16'sd-13;
        fc1_weights[28][170] = 16'sd-9;
        fc1_weights[28][171] = 16'sd-1;
        fc1_weights[28][172] = 16'sd-31;
        fc1_weights[28][173] = 16'sd-49;
        fc1_weights[28][174] = 16'sd-4;
        fc1_weights[28][175] = 16'sd18;
        fc1_weights[28][176] = 16'sd18;
        fc1_weights[28][177] = 16'sd-24;
        fc1_weights[28][178] = 16'sd15;
        fc1_weights[28][179] = 16'sd-20;
        fc1_weights[28][180] = 16'sd10;
        fc1_weights[28][181] = 16'sd-44;
        fc1_weights[28][182] = 16'sd-60;
        fc1_weights[28][183] = 16'sd-57;
        fc1_weights[28][184] = 16'sd-17;
        fc1_weights[28][185] = 16'sd-53;
        fc1_weights[28][186] = 16'sd-24;
        fc1_weights[28][187] = 16'sd50;
        fc1_weights[28][188] = 16'sd56;
        fc1_weights[28][189] = 16'sd59;
        fc1_weights[28][190] = 16'sd50;
        fc1_weights[28][191] = 16'sd11;
        fc1_weights[28][192] = 16'sd35;
        fc1_weights[28][193] = 16'sd4;
        fc1_weights[28][194] = 16'sd-11;
        fc1_weights[28][195] = 16'sd-10;
        fc1_weights[28][196] = 16'sd-2;
        fc1_weights[28][197] = 16'sd-7;
        fc1_weights[28][198] = 16'sd17;
        fc1_weights[28][199] = 16'sd-19;
        fc1_weights[28][200] = 16'sd-23;
        fc1_weights[28][201] = 16'sd11;
        fc1_weights[28][202] = 16'sd-21;
        fc1_weights[28][203] = 16'sd-2;
        fc1_weights[28][204] = 16'sd12;
        fc1_weights[28][205] = 16'sd-42;
        fc1_weights[28][206] = 16'sd-12;
        fc1_weights[28][207] = 16'sd7;
        fc1_weights[29][0] = 16'sd-68;
        fc1_weights[29][1] = 16'sd-66;
        fc1_weights[29][2] = 16'sd-12;
        fc1_weights[29][3] = 16'sd-43;
        fc1_weights[29][4] = 16'sd11;
        fc1_weights[29][5] = 16'sd0;
        fc1_weights[29][6] = 16'sd36;
        fc1_weights[29][7] = 16'sd15;
        fc1_weights[29][8] = 16'sd29;
        fc1_weights[29][9] = 16'sd40;
        fc1_weights[29][10] = 16'sd28;
        fc1_weights[29][11] = 16'sd24;
        fc1_weights[29][12] = 16'sd33;
        fc1_weights[29][13] = 16'sd13;
        fc1_weights[29][14] = 16'sd14;
        fc1_weights[29][15] = 16'sd0;
        fc1_weights[29][16] = 16'sd-52;
        fc1_weights[29][17] = 16'sd-10;
        fc1_weights[29][18] = 16'sd-10;
        fc1_weights[29][19] = 16'sd-19;
        fc1_weights[29][20] = 16'sd11;
        fc1_weights[29][21] = 16'sd15;
        fc1_weights[29][22] = 16'sd34;
        fc1_weights[29][23] = 16'sd51;
        fc1_weights[29][24] = 16'sd56;
        fc1_weights[29][25] = 16'sd60;
        fc1_weights[29][26] = 16'sd-33;
        fc1_weights[29][27] = 16'sd-59;
        fc1_weights[29][28] = 16'sd-38;
        fc1_weights[29][29] = 16'sd-22;
        fc1_weights[29][30] = 16'sd-24;
        fc1_weights[29][31] = 16'sd-9;
        fc1_weights[29][32] = 16'sd9;
        fc1_weights[29][33] = 16'sd21;
        fc1_weights[29][34] = 16'sd18;
        fc1_weights[29][35] = 16'sd39;
        fc1_weights[29][36] = 16'sd17;
        fc1_weights[29][37] = 16'sd35;
        fc1_weights[29][38] = 16'sd2;
        fc1_weights[29][39] = 16'sd-9;
        fc1_weights[29][40] = 16'sd3;
        fc1_weights[29][41] = 16'sd-25;
        fc1_weights[29][42] = 16'sd-12;
        fc1_weights[29][43] = 16'sd-53;
        fc1_weights[29][44] = 16'sd-1;
        fc1_weights[29][45] = 16'sd21;
        fc1_weights[29][46] = 16'sd30;
        fc1_weights[29][47] = 16'sd49;
        fc1_weights[29][48] = 16'sd-7;
        fc1_weights[29][49] = 16'sd41;
        fc1_weights[29][50] = 16'sd21;
        fc1_weights[29][51] = 16'sd18;
        fc1_weights[29][52] = 16'sd9;
        fc1_weights[29][53] = 16'sd-26;
        fc1_weights[29][54] = 16'sd-37;
        fc1_weights[29][55] = 16'sd-32;
        fc1_weights[29][56] = 16'sd12;
        fc1_weights[29][57] = 16'sd-8;
        fc1_weights[29][58] = 16'sd-20;
        fc1_weights[29][59] = 16'sd10;
        fc1_weights[29][60] = 16'sd16;
        fc1_weights[29][61] = 16'sd2;
        fc1_weights[29][62] = 16'sd23;
        fc1_weights[29][63] = 16'sd36;
        fc1_weights[29][64] = 16'sd12;
        fc1_weights[29][65] = 16'sd-20;
        fc1_weights[29][66] = 16'sd6;
        fc1_weights[29][67] = 16'sd-35;
        fc1_weights[29][68] = 16'sd-48;
        fc1_weights[29][69] = 16'sd28;
        fc1_weights[29][70] = 16'sd5;
        fc1_weights[29][71] = 16'sd9;
        fc1_weights[29][72] = 16'sd41;
        fc1_weights[29][73] = 16'sd39;
        fc1_weights[29][74] = 16'sd51;
        fc1_weights[29][75] = 16'sd36;
        fc1_weights[29][76] = 16'sd-12;
        fc1_weights[29][77] = 16'sd13;
        fc1_weights[29][78] = 16'sd-40;
        fc1_weights[29][79] = 16'sd30;
        fc1_weights[29][80] = 16'sd-34;
        fc1_weights[29][81] = 16'sd-35;
        fc1_weights[29][82] = 16'sd-9;
        fc1_weights[29][83] = 16'sd20;
        fc1_weights[29][84] = 16'sd-9;
        fc1_weights[29][85] = 16'sd32;
        fc1_weights[29][86] = 16'sd8;
        fc1_weights[29][87] = 16'sd47;
        fc1_weights[29][88] = 16'sd22;
        fc1_weights[29][89] = 16'sd18;
        fc1_weights[29][90] = 16'sd-5;
        fc1_weights[29][91] = 16'sd15;
        fc1_weights[29][92] = 16'sd19;
        fc1_weights[29][93] = 16'sd-33;
        fc1_weights[29][94] = 16'sd-23;
        fc1_weights[29][95] = 16'sd0;
        fc1_weights[29][96] = 16'sd-20;
        fc1_weights[29][97] = 16'sd-55;
        fc1_weights[29][98] = 16'sd3;
        fc1_weights[29][99] = 16'sd-9;
        fc1_weights[29][100] = 16'sd3;
        fc1_weights[29][101] = 16'sd12;
        fc1_weights[29][102] = 16'sd-9;
        fc1_weights[29][103] = 16'sd-3;
        fc1_weights[29][104] = 16'sd22;
        fc1_weights[29][105] = 16'sd11;
        fc1_weights[29][106] = 16'sd32;
        fc1_weights[29][107] = 16'sd-42;
        fc1_weights[29][108] = 16'sd-26;
        fc1_weights[29][109] = 16'sd-23;
        fc1_weights[29][110] = 16'sd9;
        fc1_weights[29][111] = 16'sd40;
        fc1_weights[29][112] = 16'sd-12;
        fc1_weights[29][113] = 16'sd-38;
        fc1_weights[29][114] = 16'sd4;
        fc1_weights[29][115] = 16'sd66;
        fc1_weights[29][116] = 16'sd55;
        fc1_weights[29][117] = 16'sd4;
        fc1_weights[29][118] = 16'sd-21;
        fc1_weights[29][119] = 16'sd-34;
        fc1_weights[29][120] = 16'sd-5;
        fc1_weights[29][121] = 16'sd0;
        fc1_weights[29][122] = 16'sd-14;
        fc1_weights[29][123] = 16'sd-27;
        fc1_weights[29][124] = 16'sd-18;
        fc1_weights[29][125] = 16'sd-21;
        fc1_weights[29][126] = 16'sd9;
        fc1_weights[29][127] = 16'sd-38;
        fc1_weights[29][128] = 16'sd-18;
        fc1_weights[29][129] = 16'sd8;
        fc1_weights[29][130] = 16'sd-3;
        fc1_weights[29][131] = 16'sd35;
        fc1_weights[29][132] = 16'sd13;
        fc1_weights[29][133] = 16'sd-52;
        fc1_weights[29][134] = 16'sd-49;
        fc1_weights[29][135] = 16'sd-35;
        fc1_weights[29][136] = 16'sd-15;
        fc1_weights[29][137] = 16'sd-2;
        fc1_weights[29][138] = 16'sd-16;
        fc1_weights[29][139] = 16'sd8;
        fc1_weights[29][140] = 16'sd-7;
        fc1_weights[29][141] = 16'sd78;
        fc1_weights[29][142] = 16'sd1;
        fc1_weights[29][143] = 16'sd-14;
        fc1_weights[29][144] = 16'sd-15;
        fc1_weights[29][145] = 16'sd1;
        fc1_weights[29][146] = 16'sd-19;
        fc1_weights[29][147] = 16'sd-29;
        fc1_weights[29][148] = 16'sd-55;
        fc1_weights[29][149] = 16'sd-78;
        fc1_weights[29][150] = 16'sd-17;
        fc1_weights[29][151] = 16'sd-7;
        fc1_weights[29][152] = 16'sd-16;
        fc1_weights[29][153] = 16'sd-6;
        fc1_weights[29][154] = 16'sd1;
        fc1_weights[29][155] = 16'sd10;
        fc1_weights[29][156] = 16'sd-3;
        fc1_weights[29][157] = 16'sd-14;
        fc1_weights[29][158] = 16'sd-11;
        fc1_weights[29][159] = 16'sd23;
        fc1_weights[29][160] = 16'sd15;
        fc1_weights[29][161] = 16'sd28;
        fc1_weights[29][162] = 16'sd-24;
        fc1_weights[29][163] = 16'sd-32;
        fc1_weights[29][164] = 16'sd-42;
        fc1_weights[29][165] = 16'sd-57;
        fc1_weights[29][166] = 16'sd-4;
        fc1_weights[29][167] = 16'sd-6;
        fc1_weights[29][168] = 16'sd-12;
        fc1_weights[29][169] = 16'sd-15;
        fc1_weights[29][170] = 16'sd-2;
        fc1_weights[29][171] = 16'sd26;
        fc1_weights[29][172] = 16'sd21;
        fc1_weights[29][173] = 16'sd36;
        fc1_weights[29][174] = 16'sd27;
        fc1_weights[29][175] = 16'sd-4;
        fc1_weights[29][176] = 16'sd-34;
        fc1_weights[29][177] = 16'sd-25;
        fc1_weights[29][178] = 16'sd-14;
        fc1_weights[29][179] = 16'sd-16;
        fc1_weights[29][180] = 16'sd-33;
        fc1_weights[29][181] = 16'sd-1;
        fc1_weights[29][182] = 16'sd0;
        fc1_weights[29][183] = 16'sd-15;
        fc1_weights[29][184] = 16'sd-21;
        fc1_weights[29][185] = 16'sd-29;
        fc1_weights[29][186] = 16'sd-38;
        fc1_weights[29][187] = 16'sd-40;
        fc1_weights[29][188] = 16'sd-15;
        fc1_weights[29][189] = 16'sd-12;
        fc1_weights[29][190] = 16'sd6;
        fc1_weights[29][191] = 16'sd10;
        fc1_weights[29][192] = 16'sd47;
        fc1_weights[29][193] = 16'sd13;
        fc1_weights[29][194] = 16'sd5;
        fc1_weights[29][195] = 16'sd2;
        fc1_weights[29][196] = 16'sd-4;
        fc1_weights[29][197] = 16'sd-47;
        fc1_weights[29][198] = 16'sd4;
        fc1_weights[29][199] = 16'sd27;
        fc1_weights[29][200] = 16'sd26;
        fc1_weights[29][201] = 16'sd17;
        fc1_weights[29][202] = 16'sd-12;
        fc1_weights[29][203] = 16'sd-9;
        fc1_weights[29][204] = 16'sd-16;
        fc1_weights[29][205] = 16'sd-27;
        fc1_weights[29][206] = 16'sd-20;
        fc1_weights[29][207] = 16'sd-17;
        fc1_weights[30][0] = 16'sd20;
        fc1_weights[30][1] = 16'sd48;
        fc1_weights[30][2] = 16'sd39;
        fc1_weights[30][3] = 16'sd22;
        fc1_weights[30][4] = 16'sd-8;
        fc1_weights[30][5] = 16'sd6;
        fc1_weights[30][6] = 16'sd10;
        fc1_weights[30][7] = 16'sd-2;
        fc1_weights[30][8] = 16'sd0;
        fc1_weights[30][9] = 16'sd3;
        fc1_weights[30][10] = 16'sd-18;
        fc1_weights[30][11] = 16'sd-4;
        fc1_weights[30][12] = 16'sd-54;
        fc1_weights[30][13] = 16'sd-26;
        fc1_weights[30][14] = 16'sd-28;
        fc1_weights[30][15] = 16'sd-39;
        fc1_weights[30][16] = 16'sd-8;
        fc1_weights[30][17] = 16'sd-19;
        fc1_weights[30][18] = 16'sd-30;
        fc1_weights[30][19] = 16'sd-9;
        fc1_weights[30][20] = 16'sd20;
        fc1_weights[30][21] = 16'sd-12;
        fc1_weights[30][22] = 16'sd-15;
        fc1_weights[30][23] = 16'sd2;
        fc1_weights[30][24] = 16'sd5;
        fc1_weights[30][25] = 16'sd2;
        fc1_weights[30][26] = 16'sd12;
        fc1_weights[30][27] = 16'sd13;
        fc1_weights[30][28] = 16'sd41;
        fc1_weights[30][29] = 16'sd28;
        fc1_weights[30][30] = 16'sd10;
        fc1_weights[30][31] = 16'sd18;
        fc1_weights[30][32] = 16'sd20;
        fc1_weights[30][33] = 16'sd22;
        fc1_weights[30][34] = 16'sd0;
        fc1_weights[30][35] = 16'sd10;
        fc1_weights[30][36] = 16'sd23;
        fc1_weights[30][37] = 16'sd26;
        fc1_weights[30][38] = 16'sd-3;
        fc1_weights[30][39] = 16'sd12;
        fc1_weights[30][40] = 16'sd-26;
        fc1_weights[30][41] = 16'sd-29;
        fc1_weights[30][42] = 16'sd-7;
        fc1_weights[30][43] = 16'sd-8;
        fc1_weights[30][44] = 16'sd-25;
        fc1_weights[30][45] = 16'sd-29;
        fc1_weights[30][46] = 16'sd-4;
        fc1_weights[30][47] = 16'sd18;
        fc1_weights[30][48] = 16'sd0;
        fc1_weights[30][49] = 16'sd-1;
        fc1_weights[30][50] = 16'sd3;
        fc1_weights[30][51] = 16'sd-10;
        fc1_weights[30][52] = 16'sd41;
        fc1_weights[30][53] = 16'sd22;
        fc1_weights[30][54] = 16'sd33;
        fc1_weights[30][55] = 16'sd12;
        fc1_weights[30][56] = 16'sd10;
        fc1_weights[30][57] = 16'sd25;
        fc1_weights[30][58] = 16'sd29;
        fc1_weights[30][59] = 16'sd6;
        fc1_weights[30][60] = 16'sd-18;
        fc1_weights[30][61] = 16'sd44;
        fc1_weights[30][62] = 16'sd-2;
        fc1_weights[30][63] = 16'sd15;
        fc1_weights[30][64] = 16'sd16;
        fc1_weights[30][65] = 16'sd9;
        fc1_weights[30][66] = 16'sd-33;
        fc1_weights[30][67] = 16'sd-25;
        fc1_weights[30][68] = 16'sd-8;
        fc1_weights[30][69] = 16'sd-12;
        fc1_weights[30][70] = 16'sd-31;
        fc1_weights[30][71] = 16'sd-7;
        fc1_weights[30][72] = 16'sd24;
        fc1_weights[30][73] = 16'sd23;
        fc1_weights[30][74] = 16'sd17;
        fc1_weights[30][75] = 16'sd19;
        fc1_weights[30][76] = 16'sd-3;
        fc1_weights[30][77] = 16'sd-13;
        fc1_weights[30][78] = 16'sd-2;
        fc1_weights[30][79] = 16'sd-24;
        fc1_weights[30][80] = 16'sd37;
        fc1_weights[30][81] = 16'sd-4;
        fc1_weights[30][82] = 16'sd2;
        fc1_weights[30][83] = 16'sd4;
        fc1_weights[30][84] = 16'sd28;
        fc1_weights[30][85] = 16'sd39;
        fc1_weights[30][86] = 16'sd37;
        fc1_weights[30][87] = 16'sd19;
        fc1_weights[30][88] = 16'sd0;
        fc1_weights[30][89] = 16'sd13;
        fc1_weights[30][90] = 16'sd7;
        fc1_weights[30][91] = 16'sd-15;
        fc1_weights[30][92] = 16'sd-15;
        fc1_weights[30][93] = 16'sd-14;
        fc1_weights[30][94] = 16'sd30;
        fc1_weights[30][95] = 16'sd-10;
        fc1_weights[30][96] = 16'sd-4;
        fc1_weights[30][97] = 16'sd-1;
        fc1_weights[30][98] = 16'sd7;
        fc1_weights[30][99] = 16'sd38;
        fc1_weights[30][100] = 16'sd12;
        fc1_weights[30][101] = 16'sd22;
        fc1_weights[30][102] = 16'sd11;
        fc1_weights[30][103] = 16'sd-7;
        fc1_weights[30][104] = 16'sd-25;
        fc1_weights[30][105] = 16'sd-18;
        fc1_weights[30][106] = 16'sd14;
        fc1_weights[30][107] = 16'sd12;
        fc1_weights[30][108] = 16'sd10;
        fc1_weights[30][109] = 16'sd0;
        fc1_weights[30][110] = 16'sd10;
        fc1_weights[30][111] = 16'sd-4;
        fc1_weights[30][112] = 16'sd-16;
        fc1_weights[30][113] = 16'sd-17;
        fc1_weights[30][114] = 16'sd-45;
        fc1_weights[30][115] = 16'sd-47;
        fc1_weights[30][116] = 16'sd-14;
        fc1_weights[30][117] = 16'sd-50;
        fc1_weights[30][118] = 16'sd-4;
        fc1_weights[30][119] = 16'sd12;
        fc1_weights[30][120] = 16'sd23;
        fc1_weights[30][121] = 16'sd0;
        fc1_weights[30][122] = 16'sd12;
        fc1_weights[30][123] = 16'sd5;
        fc1_weights[30][124] = 16'sd14;
        fc1_weights[30][125] = 16'sd27;
        fc1_weights[30][126] = 16'sd17;
        fc1_weights[30][127] = 16'sd20;
        fc1_weights[30][128] = 16'sd0;
        fc1_weights[30][129] = 16'sd8;
        fc1_weights[30][130] = 16'sd12;
        fc1_weights[30][131] = 16'sd24;
        fc1_weights[30][132] = 16'sd43;
        fc1_weights[30][133] = 16'sd-4;
        fc1_weights[30][134] = 16'sd0;
        fc1_weights[30][135] = 16'sd-22;
        fc1_weights[30][136] = 16'sd-23;
        fc1_weights[30][137] = 16'sd-13;
        fc1_weights[30][138] = 16'sd-47;
        fc1_weights[30][139] = 16'sd33;
        fc1_weights[30][140] = 16'sd-12;
        fc1_weights[30][141] = 16'sd-19;
        fc1_weights[30][142] = 16'sd1;
        fc1_weights[30][143] = 16'sd3;
        fc1_weights[30][144] = 16'sd-47;
        fc1_weights[30][145] = 16'sd-10;
        fc1_weights[30][146] = 16'sd14;
        fc1_weights[30][147] = 16'sd8;
        fc1_weights[30][148] = 16'sd-16;
        fc1_weights[30][149] = 16'sd24;
        fc1_weights[30][150] = 16'sd25;
        fc1_weights[30][151] = 16'sd18;
        fc1_weights[30][152] = 16'sd28;
        fc1_weights[30][153] = 16'sd17;
        fc1_weights[30][154] = 16'sd19;
        fc1_weights[30][155] = 16'sd23;
        fc1_weights[30][156] = 16'sd5;
        fc1_weights[30][157] = 16'sd-26;
        fc1_weights[30][158] = 16'sd3;
        fc1_weights[30][159] = 16'sd-19;
        fc1_weights[30][160] = 16'sd16;
        fc1_weights[30][161] = 16'sd13;
        fc1_weights[30][162] = 16'sd-13;
        fc1_weights[30][163] = 16'sd21;
        fc1_weights[30][164] = 16'sd33;
        fc1_weights[30][165] = 16'sd30;
        fc1_weights[30][166] = 16'sd0;
        fc1_weights[30][167] = 16'sd17;
        fc1_weights[30][168] = 16'sd-16;
        fc1_weights[30][169] = 16'sd4;
        fc1_weights[30][170] = 16'sd-2;
        fc1_weights[30][171] = 16'sd-57;
        fc1_weights[30][172] = 16'sd-16;
        fc1_weights[30][173] = 16'sd1;
        fc1_weights[30][174] = 16'sd-6;
        fc1_weights[30][175] = 16'sd-12;
        fc1_weights[30][176] = 16'sd46;
        fc1_weights[30][177] = 16'sd-8;
        fc1_weights[30][178] = 16'sd45;
        fc1_weights[30][179] = 16'sd37;
        fc1_weights[30][180] = 16'sd-9;
        fc1_weights[30][181] = 16'sd12;
        fc1_weights[30][182] = 16'sd-8;
        fc1_weights[30][183] = 16'sd-2;
        fc1_weights[30][184] = 16'sd5;
        fc1_weights[30][185] = 16'sd-8;
        fc1_weights[30][186] = 16'sd-19;
        fc1_weights[30][187] = 16'sd5;
        fc1_weights[30][188] = 16'sd7;
        fc1_weights[30][189] = 16'sd16;
        fc1_weights[30][190] = 16'sd0;
        fc1_weights[30][191] = 16'sd21;
        fc1_weights[30][192] = 16'sd32;
        fc1_weights[30][193] = 16'sd20;
        fc1_weights[30][194] = 16'sd-32;
        fc1_weights[30][195] = 16'sd-12;
        fc1_weights[30][196] = 16'sd7;
        fc1_weights[30][197] = 16'sd-4;
        fc1_weights[30][198] = 16'sd-20;
        fc1_weights[30][199] = 16'sd0;
        fc1_weights[30][200] = 16'sd20;
        fc1_weights[30][201] = 16'sd7;
        fc1_weights[30][202] = 16'sd-25;
        fc1_weights[30][203] = 16'sd17;
        fc1_weights[30][204] = 16'sd19;
        fc1_weights[30][205] = 16'sd8;
        fc1_weights[30][206] = 16'sd-5;
        fc1_weights[30][207] = 16'sd16;
        fc1_weights[31][0] = 16'sd5;
        fc1_weights[31][1] = 16'sd-1;
        fc1_weights[31][2] = 16'sd-10;
        fc1_weights[31][3] = 16'sd9;
        fc1_weights[31][4] = 16'sd-9;
        fc1_weights[31][5] = 16'sd8;
        fc1_weights[31][6] = 16'sd-5;
        fc1_weights[31][7] = 16'sd-20;
        fc1_weights[31][8] = 16'sd-6;
        fc1_weights[31][9] = 16'sd-16;
        fc1_weights[31][10] = 16'sd-53;
        fc1_weights[31][11] = 16'sd-49;
        fc1_weights[31][12] = 16'sd69;
        fc1_weights[31][13] = 16'sd91;
        fc1_weights[31][14] = 16'sd102;
        fc1_weights[31][15] = 16'sd26;
        fc1_weights[31][16] = 16'sd12;
        fc1_weights[31][17] = 16'sd0;
        fc1_weights[31][18] = 16'sd-11;
        fc1_weights[31][19] = 16'sd6;
        fc1_weights[31][20] = 16'sd-11;
        fc1_weights[31][21] = 16'sd7;
        fc1_weights[31][22] = 16'sd-13;
        fc1_weights[31][23] = 16'sd42;
        fc1_weights[31][24] = 16'sd-22;
        fc1_weights[31][25] = 16'sd-14;
        fc1_weights[31][26] = 16'sd-28;
        fc1_weights[31][27] = 16'sd-16;
        fc1_weights[31][28] = 16'sd31;
        fc1_weights[31][29] = 16'sd-22;
        fc1_weights[31][30] = 16'sd-15;
        fc1_weights[31][31] = 16'sd3;
        fc1_weights[31][32] = 16'sd-8;
        fc1_weights[31][33] = 16'sd48;
        fc1_weights[31][34] = 16'sd-24;
        fc1_weights[31][35] = 16'sd11;
        fc1_weights[31][36] = 16'sd-34;
        fc1_weights[31][37] = 16'sd-46;
        fc1_weights[31][38] = 16'sd-10;
        fc1_weights[31][39] = 16'sd44;
        fc1_weights[31][40] = 16'sd-24;
        fc1_weights[31][41] = 16'sd60;
        fc1_weights[31][42] = 16'sd43;
        fc1_weights[31][43] = 16'sd-10;
        fc1_weights[31][44] = 16'sd-21;
        fc1_weights[31][45] = 16'sd-10;
        fc1_weights[31][46] = 16'sd-20;
        fc1_weights[31][47] = 16'sd19;
        fc1_weights[31][48] = 16'sd-36;
        fc1_weights[31][49] = 16'sd-40;
        fc1_weights[31][50] = 16'sd-23;
        fc1_weights[31][51] = 16'sd-32;
        fc1_weights[31][52] = 16'sd22;
        fc1_weights[31][53] = 16'sd-37;
        fc1_weights[31][54] = 16'sd31;
        fc1_weights[31][55] = 16'sd55;
        fc1_weights[31][56] = 16'sd11;
        fc1_weights[31][57] = 16'sd2;
        fc1_weights[31][58] = 16'sd-17;
        fc1_weights[31][59] = 16'sd-14;
        fc1_weights[31][60] = 16'sd-13;
        fc1_weights[31][61] = 16'sd-7;
        fc1_weights[31][62] = 16'sd16;
        fc1_weights[31][63] = 16'sd-7;
        fc1_weights[31][64] = 16'sd-16;
        fc1_weights[31][65] = 16'sd17;
        fc1_weights[31][66] = 16'sd10;
        fc1_weights[31][67] = 16'sd50;
        fc1_weights[31][68] = 16'sd-52;
        fc1_weights[31][69] = 16'sd11;
        fc1_weights[31][70] = 16'sd15;
        fc1_weights[31][71] = 16'sd-13;
        fc1_weights[31][72] = 16'sd-63;
        fc1_weights[31][73] = 16'sd40;
        fc1_weights[31][74] = 16'sd16;
        fc1_weights[31][75] = 16'sd1;
        fc1_weights[31][76] = 16'sd-45;
        fc1_weights[31][77] = 16'sd-42;
        fc1_weights[31][78] = 16'sd-7;
        fc1_weights[31][79] = 16'sd-28;
        fc1_weights[31][80] = 16'sd-7;
        fc1_weights[31][81] = 16'sd77;
        fc1_weights[31][82] = 16'sd60;
        fc1_weights[31][83] = 16'sd104;
        fc1_weights[31][84] = 16'sd60;
        fc1_weights[31][85] = 16'sd39;
        fc1_weights[31][86] = 16'sd53;
        fc1_weights[31][87] = 16'sd1;
        fc1_weights[31][88] = 16'sd41;
        fc1_weights[31][89] = 16'sd-50;
        fc1_weights[31][90] = 16'sd-141;
        fc1_weights[31][91] = 16'sd-40;
        fc1_weights[31][92] = 16'sd-26;
        fc1_weights[31][93] = 16'sd25;
        fc1_weights[31][94] = 16'sd-22;
        fc1_weights[31][95] = 16'sd36;
        fc1_weights[31][96] = 16'sd51;
        fc1_weights[31][97] = 16'sd-19;
        fc1_weights[31][98] = 16'sd-6;
        fc1_weights[31][99] = 16'sd32;
        fc1_weights[31][100] = 16'sd5;
        fc1_weights[31][101] = 16'sd18;
        fc1_weights[31][102] = 16'sd-3;
        fc1_weights[31][103] = 16'sd10;
        fc1_weights[31][104] = 16'sd12;
        fc1_weights[31][105] = 16'sd-35;
        fc1_weights[31][106] = 16'sd27;
        fc1_weights[31][107] = 16'sd13;
        fc1_weights[31][108] = 16'sd-6;
        fc1_weights[31][109] = 16'sd-4;
        fc1_weights[31][110] = 16'sd-18;
        fc1_weights[31][111] = 16'sd6;
        fc1_weights[31][112] = 16'sd29;
        fc1_weights[31][113] = 16'sd-12;
        fc1_weights[31][114] = 16'sd17;
        fc1_weights[31][115] = 16'sd-15;
        fc1_weights[31][116] = 16'sd70;
        fc1_weights[31][117] = 16'sd-7;
        fc1_weights[31][118] = 16'sd-6;
        fc1_weights[31][119] = 16'sd22;
        fc1_weights[31][120] = 16'sd48;
        fc1_weights[31][121] = 16'sd28;
        fc1_weights[31][122] = 16'sd24;
        fc1_weights[31][123] = 16'sd4;
        fc1_weights[31][124] = 16'sd17;
        fc1_weights[31][125] = 16'sd44;
        fc1_weights[31][126] = 16'sd40;
        fc1_weights[31][127] = 16'sd-25;
        fc1_weights[31][128] = 16'sd-26;
        fc1_weights[31][129] = 16'sd32;
        fc1_weights[31][130] = 16'sd47;
        fc1_weights[31][131] = 16'sd-2;
        fc1_weights[31][132] = 16'sd-1;
        fc1_weights[31][133] = 16'sd-37;
        fc1_weights[31][134] = 16'sd-29;
        fc1_weights[31][135] = 16'sd-10;
        fc1_weights[31][136] = 16'sd-22;
        fc1_weights[31][137] = 16'sd1;
        fc1_weights[31][138] = 16'sd-36;
        fc1_weights[31][139] = 16'sd14;
        fc1_weights[31][140] = 16'sd-41;
        fc1_weights[31][141] = 16'sd-8;
        fc1_weights[31][142] = 16'sd-70;
        fc1_weights[31][143] = 16'sd12;
        fc1_weights[31][144] = 16'sd-5;
        fc1_weights[31][145] = 16'sd31;
        fc1_weights[31][146] = 16'sd36;
        fc1_weights[31][147] = 16'sd39;
        fc1_weights[31][148] = 16'sd4;
        fc1_weights[31][149] = 16'sd38;
        fc1_weights[31][150] = 16'sd25;
        fc1_weights[31][151] = 16'sd71;
        fc1_weights[31][152] = 16'sd-4;
        fc1_weights[31][153] = 16'sd-14;
        fc1_weights[31][154] = 16'sd19;
        fc1_weights[31][155] = 16'sd-40;
        fc1_weights[31][156] = 16'sd-25;
        fc1_weights[31][157] = 16'sd-25;
        fc1_weights[31][158] = 16'sd9;
        fc1_weights[31][159] = 16'sd0;
        fc1_weights[31][160] = 16'sd8;
        fc1_weights[31][161] = 16'sd43;
        fc1_weights[31][162] = 16'sd-70;
        fc1_weights[31][163] = 16'sd-33;
        fc1_weights[31][164] = 16'sd-37;
        fc1_weights[31][165] = 16'sd-66;
        fc1_weights[31][166] = 16'sd-93;
        fc1_weights[31][167] = 16'sd-52;
        fc1_weights[31][168] = 16'sd-23;
        fc1_weights[31][169] = 16'sd10;
        fc1_weights[31][170] = 16'sd-19;
        fc1_weights[31][171] = 16'sd-45;
        fc1_weights[31][172] = 16'sd-20;
        fc1_weights[31][173] = 16'sd0;
        fc1_weights[31][174] = 16'sd21;
        fc1_weights[31][175] = 16'sd-11;
        fc1_weights[31][176] = 16'sd30;
        fc1_weights[31][177] = 16'sd-39;
        fc1_weights[31][178] = 16'sd58;
        fc1_weights[31][179] = 16'sd-19;
        fc1_weights[31][180] = 16'sd49;
        fc1_weights[31][181] = 16'sd-3;
        fc1_weights[31][182] = 16'sd2;
        fc1_weights[31][183] = 16'sd-7;
        fc1_weights[31][184] = 16'sd34;
        fc1_weights[31][185] = 16'sd1;
        fc1_weights[31][186] = 16'sd6;
        fc1_weights[31][187] = 16'sd11;
        fc1_weights[31][188] = 16'sd-15;
        fc1_weights[31][189] = 16'sd15;
        fc1_weights[31][190] = 16'sd-2;
        fc1_weights[31][191] = 16'sd-66;
        fc1_weights[31][192] = 16'sd0;
        fc1_weights[31][193] = 16'sd-24;
        fc1_weights[31][194] = 16'sd-35;
        fc1_weights[31][195] = 16'sd-24;
        fc1_weights[31][196] = 16'sd8;
        fc1_weights[31][197] = 16'sd-65;
        fc1_weights[31][198] = 16'sd-11;
        fc1_weights[31][199] = 16'sd0;
        fc1_weights[31][200] = 16'sd7;
        fc1_weights[31][201] = 16'sd14;
        fc1_weights[31][202] = 16'sd-26;
        fc1_weights[31][203] = 16'sd-24;
        fc1_weights[31][204] = 16'sd-3;
        fc1_weights[31][205] = 16'sd-17;
        fc1_weights[31][206] = 16'sd18;
        fc1_weights[31][207] = 16'sd34;
        fc1_weights[32][0] = 16'sd2;
        fc1_weights[32][1] = 16'sd-31;
        fc1_weights[32][2] = 16'sd-94;
        fc1_weights[32][3] = 16'sd-60;
        fc1_weights[32][4] = 16'sd27;
        fc1_weights[32][5] = 16'sd-57;
        fc1_weights[32][6] = 16'sd29;
        fc1_weights[32][7] = 16'sd-38;
        fc1_weights[32][8] = 16'sd64;
        fc1_weights[32][9] = 16'sd17;
        fc1_weights[32][10] = 16'sd5;
        fc1_weights[32][11] = 16'sd40;
        fc1_weights[32][12] = 16'sd93;
        fc1_weights[32][13] = 16'sd10;
        fc1_weights[32][14] = 16'sd-16;
        fc1_weights[32][15] = 16'sd-8;
        fc1_weights[32][16] = 16'sd73;
        fc1_weights[32][17] = 16'sd0;
        fc1_weights[32][18] = 16'sd0;
        fc1_weights[32][19] = 16'sd-25;
        fc1_weights[32][20] = 16'sd-27;
        fc1_weights[32][21] = 16'sd2;
        fc1_weights[32][22] = 16'sd45;
        fc1_weights[32][23] = 16'sd22;
        fc1_weights[32][24] = 16'sd-16;
        fc1_weights[32][25] = 16'sd16;
        fc1_weights[32][26] = 16'sd18;
        fc1_weights[32][27] = 16'sd-21;
        fc1_weights[32][28] = 16'sd-68;
        fc1_weights[32][29] = 16'sd-84;
        fc1_weights[32][30] = 16'sd-40;
        fc1_weights[32][31] = 16'sd-51;
        fc1_weights[32][32] = 16'sd17;
        fc1_weights[32][33] = 16'sd87;
        fc1_weights[32][34] = 16'sd-16;
        fc1_weights[32][35] = 16'sd-23;
        fc1_weights[32][36] = 16'sd-16;
        fc1_weights[32][37] = 16'sd-3;
        fc1_weights[32][38] = 16'sd66;
        fc1_weights[32][39] = 16'sd-20;
        fc1_weights[32][40] = 16'sd-80;
        fc1_weights[32][41] = 16'sd-26;
        fc1_weights[32][42] = 16'sd64;
        fc1_weights[32][43] = 16'sd20;
        fc1_weights[32][44] = 16'sd46;
        fc1_weights[32][45] = 16'sd10;
        fc1_weights[32][46] = 16'sd94;
        fc1_weights[32][47] = 16'sd22;
        fc1_weights[32][48] = 16'sd23;
        fc1_weights[32][49] = 16'sd-46;
        fc1_weights[32][50] = 16'sd23;
        fc1_weights[32][51] = 16'sd64;
        fc1_weights[32][52] = 16'sd-11;
        fc1_weights[32][53] = 16'sd-18;
        fc1_weights[32][54] = 16'sd15;
        fc1_weights[32][55] = 16'sd-29;
        fc1_weights[32][56] = 16'sd0;
        fc1_weights[32][57] = 16'sd-30;
        fc1_weights[32][58] = 16'sd11;
        fc1_weights[32][59] = 16'sd-33;
        fc1_weights[32][60] = 16'sd-94;
        fc1_weights[32][61] = 16'sd1;
        fc1_weights[32][62] = 16'sd49;
        fc1_weights[32][63] = 16'sd-6;
        fc1_weights[32][64] = 16'sd-52;
        fc1_weights[32][65] = 16'sd48;
        fc1_weights[32][66] = 16'sd19;
        fc1_weights[32][67] = 16'sd27;
        fc1_weights[32][68] = 16'sd81;
        fc1_weights[32][69] = 16'sd10;
        fc1_weights[32][70] = 16'sd-64;
        fc1_weights[32][71] = 16'sd-4;
        fc1_weights[32][72] = 16'sd-41;
        fc1_weights[32][73] = 16'sd16;
        fc1_weights[32][74] = 16'sd-6;
        fc1_weights[32][75] = 16'sd-2;
        fc1_weights[32][76] = 16'sd21;
        fc1_weights[32][77] = 16'sd1;
        fc1_weights[32][78] = 16'sd-21;
        fc1_weights[32][79] = 16'sd-35;
        fc1_weights[32][80] = 16'sd13;
        fc1_weights[32][81] = 16'sd29;
        fc1_weights[32][82] = 16'sd5;
        fc1_weights[32][83] = 16'sd-18;
        fc1_weights[32][84] = 16'sd-10;
        fc1_weights[32][85] = 16'sd4;
        fc1_weights[32][86] = 16'sd19;
        fc1_weights[32][87] = 16'sd17;
        fc1_weights[32][88] = 16'sd21;
        fc1_weights[32][89] = 16'sd48;
        fc1_weights[32][90] = 16'sd-51;
        fc1_weights[32][91] = 16'sd65;
        fc1_weights[32][92] = 16'sd38;
        fc1_weights[32][93] = 16'sd-29;
        fc1_weights[32][94] = 16'sd53;
        fc1_weights[32][95] = 16'sd22;
        fc1_weights[32][96] = 16'sd-1;
        fc1_weights[32][97] = 16'sd-39;
        fc1_weights[32][98] = 16'sd-30;
        fc1_weights[32][99] = 16'sd98;
        fc1_weights[32][100] = 16'sd50;
        fc1_weights[32][101] = 16'sd1;
        fc1_weights[32][102] = 16'sd31;
        fc1_weights[32][103] = 16'sd25;
        fc1_weights[32][104] = 16'sd-33;
        fc1_weights[32][105] = 16'sd28;
        fc1_weights[32][106] = 16'sd-6;
        fc1_weights[32][107] = 16'sd23;
        fc1_weights[32][108] = 16'sd10;
        fc1_weights[32][109] = 16'sd47;
        fc1_weights[32][110] = 16'sd-1;
        fc1_weights[32][111] = 16'sd-39;
        fc1_weights[32][112] = 16'sd-121;
        fc1_weights[32][113] = 16'sd-52;
        fc1_weights[32][114] = 16'sd-1;
        fc1_weights[32][115] = 16'sd5;
        fc1_weights[32][116] = 16'sd52;
        fc1_weights[32][117] = 16'sd24;
        fc1_weights[32][118] = 16'sd-52;
        fc1_weights[32][119] = 16'sd25;
        fc1_weights[32][120] = 16'sd77;
        fc1_weights[32][121] = 16'sd-24;
        fc1_weights[32][122] = 16'sd-53;
        fc1_weights[32][123] = 16'sd-6;
        fc1_weights[32][124] = 16'sd26;
        fc1_weights[32][125] = 16'sd46;
        fc1_weights[32][126] = 16'sd-20;
        fc1_weights[32][127] = 16'sd-28;
        fc1_weights[32][128] = 16'sd-24;
        fc1_weights[32][129] = 16'sd-30;
        fc1_weights[32][130] = 16'sd-2;
        fc1_weights[32][131] = 16'sd-23;
        fc1_weights[32][132] = 16'sd-2;
        fc1_weights[32][133] = 16'sd31;
        fc1_weights[32][134] = 16'sd47;
        fc1_weights[32][135] = 16'sd38;
        fc1_weights[32][136] = 16'sd24;
        fc1_weights[32][137] = 16'sd21;
        fc1_weights[32][138] = 16'sd-106;
        fc1_weights[32][139] = 16'sd-12;
        fc1_weights[32][140] = 16'sd5;
        fc1_weights[32][141] = 16'sd-17;
        fc1_weights[32][142] = 16'sd0;
        fc1_weights[32][143] = 16'sd-5;
        fc1_weights[32][144] = 16'sd-67;
        fc1_weights[32][145] = 16'sd9;
        fc1_weights[32][146] = 16'sd44;
        fc1_weights[32][147] = 16'sd17;
        fc1_weights[32][148] = 16'sd-11;
        fc1_weights[32][149] = 16'sd33;
        fc1_weights[32][150] = 16'sd-62;
        fc1_weights[32][151] = 16'sd-65;
        fc1_weights[32][152] = 16'sd-55;
        fc1_weights[32][153] = 16'sd-88;
        fc1_weights[32][154] = 16'sd-55;
        fc1_weights[32][155] = 16'sd-82;
        fc1_weights[32][156] = 16'sd24;
        fc1_weights[32][157] = 16'sd16;
        fc1_weights[32][158] = 16'sd22;
        fc1_weights[32][159] = 16'sd10;
        fc1_weights[32][160] = 16'sd-1;
        fc1_weights[32][161] = 16'sd50;
        fc1_weights[32][162] = 16'sd-37;
        fc1_weights[32][163] = 16'sd21;
        fc1_weights[32][164] = 16'sd-9;
        fc1_weights[32][165] = 16'sd64;
        fc1_weights[32][166] = 16'sd38;
        fc1_weights[32][167] = 16'sd33;
        fc1_weights[32][168] = 16'sd31;
        fc1_weights[32][169] = 16'sd91;
        fc1_weights[32][170] = 16'sd65;
        fc1_weights[32][171] = 16'sd86;
        fc1_weights[32][172] = 16'sd-24;
        fc1_weights[32][173] = 16'sd53;
        fc1_weights[32][174] = 16'sd81;
        fc1_weights[32][175] = 16'sd87;
        fc1_weights[32][176] = 16'sd44;
        fc1_weights[32][177] = 16'sd-22;
        fc1_weights[32][178] = 16'sd27;
        fc1_weights[32][179] = 16'sd-43;
        fc1_weights[32][180] = 16'sd-69;
        fc1_weights[32][181] = 16'sd-94;
        fc1_weights[32][182] = 16'sd24;
        fc1_weights[32][183] = 16'sd32;
        fc1_weights[32][184] = 16'sd56;
        fc1_weights[32][185] = 16'sd31;
        fc1_weights[32][186] = 16'sd6;
        fc1_weights[32][187] = 16'sd23;
        fc1_weights[32][188] = 16'sd51;
        fc1_weights[32][189] = 16'sd39;
        fc1_weights[32][190] = 16'sd-24;
        fc1_weights[32][191] = 16'sd-17;
        fc1_weights[32][192] = 16'sd-46;
        fc1_weights[32][193] = 16'sd13;
        fc1_weights[32][194] = 16'sd10;
        fc1_weights[32][195] = 16'sd61;
        fc1_weights[32][196] = 16'sd65;
        fc1_weights[32][197] = 16'sd27;
        fc1_weights[32][198] = 16'sd71;
        fc1_weights[32][199] = 16'sd12;
        fc1_weights[32][200] = 16'sd-29;
        fc1_weights[32][201] = 16'sd8;
        fc1_weights[32][202] = 16'sd9;
        fc1_weights[32][203] = 16'sd-29;
        fc1_weights[32][204] = 16'sd-79;
        fc1_weights[32][205] = 16'sd-46;
        fc1_weights[32][206] = 16'sd-92;
        fc1_weights[32][207] = 16'sd-56;
        fc1_weights[33][0] = 16'sd20;
        fc1_weights[33][1] = 16'sd5;
        fc1_weights[33][2] = 16'sd2;
        fc1_weights[33][3] = 16'sd113;
        fc1_weights[33][4] = 16'sd26;
        fc1_weights[33][5] = 16'sd32;
        fc1_weights[33][6] = 16'sd24;
        fc1_weights[33][7] = 16'sd-6;
        fc1_weights[33][8] = 16'sd13;
        fc1_weights[33][9] = 16'sd83;
        fc1_weights[33][10] = 16'sd66;
        fc1_weights[33][11] = 16'sd85;
        fc1_weights[33][12] = 16'sd115;
        fc1_weights[33][13] = 16'sd60;
        fc1_weights[33][14] = 16'sd89;
        fc1_weights[33][15] = 16'sd34;
        fc1_weights[33][16] = 16'sd32;
        fc1_weights[33][17] = 16'sd31;
        fc1_weights[33][18] = 16'sd6;
        fc1_weights[33][19] = 16'sd1;
        fc1_weights[33][20] = 16'sd-55;
        fc1_weights[33][21] = 16'sd-18;
        fc1_weights[33][22] = 16'sd17;
        fc1_weights[33][23] = 16'sd38;
        fc1_weights[33][24] = 16'sd18;
        fc1_weights[33][25] = 16'sd0;
        fc1_weights[33][26] = 16'sd0;
        fc1_weights[33][27] = 16'sd-4;
        fc1_weights[33][28] = 16'sd31;
        fc1_weights[33][29] = 16'sd-3;
        fc1_weights[33][30] = 16'sd-70;
        fc1_weights[33][31] = 16'sd-47;
        fc1_weights[33][32] = 16'sd-35;
        fc1_weights[33][33] = 16'sd43;
        fc1_weights[33][34] = 16'sd-48;
        fc1_weights[33][35] = 16'sd23;
        fc1_weights[33][36] = 16'sd34;
        fc1_weights[33][37] = 16'sd-3;
        fc1_weights[33][38] = 16'sd46;
        fc1_weights[33][39] = 16'sd24;
        fc1_weights[33][40] = 16'sd1;
        fc1_weights[33][41] = 16'sd21;
        fc1_weights[33][42] = 16'sd24;
        fc1_weights[33][43] = 16'sd14;
        fc1_weights[33][44] = 16'sd41;
        fc1_weights[33][45] = 16'sd36;
        fc1_weights[33][46] = 16'sd24;
        fc1_weights[33][47] = 16'sd1;
        fc1_weights[33][48] = 16'sd23;
        fc1_weights[33][49] = 16'sd-17;
        fc1_weights[33][50] = 16'sd24;
        fc1_weights[33][51] = 16'sd-7;
        fc1_weights[33][52] = 16'sd49;
        fc1_weights[33][53] = 16'sd48;
        fc1_weights[33][54] = 16'sd-9;
        fc1_weights[33][55] = 16'sd-23;
        fc1_weights[33][56] = 16'sd-16;
        fc1_weights[33][57] = 16'sd-19;
        fc1_weights[33][58] = 16'sd19;
        fc1_weights[33][59] = 16'sd-33;
        fc1_weights[33][60] = 16'sd-43;
        fc1_weights[33][61] = 16'sd4;
        fc1_weights[33][62] = 16'sd-11;
        fc1_weights[33][63] = 16'sd-19;
        fc1_weights[33][64] = 16'sd28;
        fc1_weights[33][65] = 16'sd58;
        fc1_weights[33][66] = 16'sd-29;
        fc1_weights[33][67] = 16'sd1;
        fc1_weights[33][68] = 16'sd47;
        fc1_weights[33][69] = 16'sd18;
        fc1_weights[33][70] = 16'sd0;
        fc1_weights[33][71] = 16'sd-4;
        fc1_weights[33][72] = 16'sd-17;
        fc1_weights[33][73] = 16'sd55;
        fc1_weights[33][74] = 16'sd-22;
        fc1_weights[33][75] = 16'sd-11;
        fc1_weights[33][76] = 16'sd-25;
        fc1_weights[33][77] = 16'sd-36;
        fc1_weights[33][78] = 16'sd-8;
        fc1_weights[33][79] = 16'sd-33;
        fc1_weights[33][80] = 16'sd-12;
        fc1_weights[33][81] = 16'sd-36;
        fc1_weights[33][82] = 16'sd38;
        fc1_weights[33][83] = 16'sd-42;
        fc1_weights[33][84] = 16'sd5;
        fc1_weights[33][85] = 16'sd1;
        fc1_weights[33][86] = 16'sd-28;
        fc1_weights[33][87] = 16'sd-73;
        fc1_weights[33][88] = 16'sd-96;
        fc1_weights[33][89] = 16'sd-74;
        fc1_weights[33][90] = 16'sd-2;
        fc1_weights[33][91] = 16'sd-41;
        fc1_weights[33][92] = 16'sd-69;
        fc1_weights[33][93] = 16'sd-26;
        fc1_weights[33][94] = 16'sd16;
        fc1_weights[33][95] = 16'sd-80;
        fc1_weights[33][96] = 16'sd62;
        fc1_weights[33][97] = 16'sd-25;
        fc1_weights[33][98] = 16'sd8;
        fc1_weights[33][99] = 16'sd-8;
        fc1_weights[33][100] = 16'sd-68;
        fc1_weights[33][101] = 16'sd-5;
        fc1_weights[33][102] = 16'sd-48;
        fc1_weights[33][103] = 16'sd-7;
        fc1_weights[33][104] = 16'sd-10;
        fc1_weights[33][105] = 16'sd57;
        fc1_weights[33][106] = 16'sd-9;
        fc1_weights[33][107] = 16'sd10;
        fc1_weights[33][108] = 16'sd2;
        fc1_weights[33][109] = 16'sd-11;
        fc1_weights[33][110] = 16'sd-10;
        fc1_weights[33][111] = 16'sd-26;
        fc1_weights[33][112] = 16'sd-101;
        fc1_weights[33][113] = 16'sd2;
        fc1_weights[33][114] = 16'sd-11;
        fc1_weights[33][115] = 16'sd37;
        fc1_weights[33][116] = 16'sd-2;
        fc1_weights[33][117] = 16'sd-83;
        fc1_weights[33][118] = 16'sd-17;
        fc1_weights[33][119] = 16'sd-69;
        fc1_weights[33][120] = 16'sd-20;
        fc1_weights[33][121] = 16'sd-42;
        fc1_weights[33][122] = 16'sd3;
        fc1_weights[33][123] = 16'sd-76;
        fc1_weights[33][124] = 16'sd-1;
        fc1_weights[33][125] = 16'sd53;
        fc1_weights[33][126] = 16'sd23;
        fc1_weights[33][127] = 16'sd-1;
        fc1_weights[33][128] = 16'sd-55;
        fc1_weights[33][129] = 16'sd-42;
        fc1_weights[33][130] = 16'sd34;
        fc1_weights[33][131] = 16'sd41;
        fc1_weights[33][132] = 16'sd-15;
        fc1_weights[33][133] = 16'sd-19;
        fc1_weights[33][134] = 16'sd26;
        fc1_weights[33][135] = 16'sd-44;
        fc1_weights[33][136] = 16'sd-44;
        fc1_weights[33][137] = 16'sd-11;
        fc1_weights[33][138] = 16'sd39;
        fc1_weights[33][139] = 16'sd44;
        fc1_weights[33][140] = 16'sd43;
        fc1_weights[33][141] = 16'sd5;
        fc1_weights[33][142] = 16'sd-41;
        fc1_weights[33][143] = 16'sd21;
        fc1_weights[33][144] = 16'sd-52;
        fc1_weights[33][145] = 16'sd50;
        fc1_weights[33][146] = 16'sd-5;
        fc1_weights[33][147] = 16'sd-34;
        fc1_weights[33][148] = 16'sd-42;
        fc1_weights[33][149] = 16'sd-17;
        fc1_weights[33][150] = 16'sd17;
        fc1_weights[33][151] = 16'sd-3;
        fc1_weights[33][152] = 16'sd44;
        fc1_weights[33][153] = 16'sd-6;
        fc1_weights[33][154] = 16'sd29;
        fc1_weights[33][155] = 16'sd-6;
        fc1_weights[33][156] = 16'sd-32;
        fc1_weights[33][157] = 16'sd-60;
        fc1_weights[33][158] = 16'sd-20;
        fc1_weights[33][159] = 16'sd-16;
        fc1_weights[33][160] = 16'sd88;
        fc1_weights[33][161] = 16'sd41;
        fc1_weights[33][162] = 16'sd-43;
        fc1_weights[33][163] = 16'sd-3;
        fc1_weights[33][164] = 16'sd29;
        fc1_weights[33][165] = 16'sd82;
        fc1_weights[33][166] = 16'sd70;
        fc1_weights[33][167] = 16'sd66;
        fc1_weights[33][168] = 16'sd38;
        fc1_weights[33][169] = 16'sd20;
        fc1_weights[33][170] = 16'sd-22;
        fc1_weights[33][171] = 16'sd-36;
        fc1_weights[33][172] = 16'sd-43;
        fc1_weights[33][173] = 16'sd-23;
        fc1_weights[33][174] = 16'sd-20;
        fc1_weights[33][175] = 16'sd30;
        fc1_weights[33][176] = 16'sd17;
        fc1_weights[33][177] = 16'sd-44;
        fc1_weights[33][178] = 16'sd49;
        fc1_weights[33][179] = 16'sd45;
        fc1_weights[33][180] = 16'sd-21;
        fc1_weights[33][181] = 16'sd-25;
        fc1_weights[33][182] = 16'sd-34;
        fc1_weights[33][183] = 16'sd-25;
        fc1_weights[33][184] = 16'sd13;
        fc1_weights[33][185] = 16'sd-22;
        fc1_weights[33][186] = 16'sd-27;
        fc1_weights[33][187] = 16'sd67;
        fc1_weights[33][188] = 16'sd67;
        fc1_weights[33][189] = 16'sd53;
        fc1_weights[33][190] = 16'sd26;
        fc1_weights[33][191] = 16'sd42;
        fc1_weights[33][192] = 16'sd59;
        fc1_weights[33][193] = 16'sd62;
        fc1_weights[33][194] = 16'sd-10;
        fc1_weights[33][195] = 16'sd9;
        fc1_weights[33][196] = 16'sd-3;
        fc1_weights[33][197] = 16'sd-80;
        fc1_weights[33][198] = 16'sd4;
        fc1_weights[33][199] = 16'sd-17;
        fc1_weights[33][200] = 16'sd-6;
        fc1_weights[33][201] = 16'sd-3;
        fc1_weights[33][202] = 16'sd-25;
        fc1_weights[33][203] = 16'sd10;
        fc1_weights[33][204] = 16'sd30;
        fc1_weights[33][205] = 16'sd5;
        fc1_weights[33][206] = 16'sd12;
        fc1_weights[33][207] = 16'sd1;
        fc1_weights[34][0] = 16'sd40;
        fc1_weights[34][1] = 16'sd-36;
        fc1_weights[34][2] = 16'sd-45;
        fc1_weights[34][3] = 16'sd24;
        fc1_weights[34][4] = 16'sd-1;
        fc1_weights[34][5] = 16'sd25;
        fc1_weights[34][6] = 16'sd10;
        fc1_weights[34][7] = 16'sd59;
        fc1_weights[34][8] = 16'sd-12;
        fc1_weights[34][9] = 16'sd-1;
        fc1_weights[34][10] = 16'sd7;
        fc1_weights[34][11] = 16'sd54;
        fc1_weights[34][12] = 16'sd35;
        fc1_weights[34][13] = 16'sd-15;
        fc1_weights[34][14] = 16'sd-63;
        fc1_weights[34][15] = 16'sd-24;
        fc1_weights[34][16] = 16'sd-35;
        fc1_weights[34][17] = 16'sd-16;
        fc1_weights[34][18] = 16'sd18;
        fc1_weights[34][19] = 16'sd5;
        fc1_weights[34][20] = 16'sd-3;
        fc1_weights[34][21] = 16'sd-17;
        fc1_weights[34][22] = 16'sd-50;
        fc1_weights[34][23] = 16'sd7;
        fc1_weights[34][24] = 16'sd31;
        fc1_weights[34][25] = 16'sd-38;
        fc1_weights[34][26] = 16'sd-21;
        fc1_weights[34][27] = 16'sd-35;
        fc1_weights[34][28] = 16'sd-70;
        fc1_weights[34][29] = 16'sd-20;
        fc1_weights[34][30] = 16'sd20;
        fc1_weights[34][31] = 16'sd35;
        fc1_weights[34][32] = 16'sd29;
        fc1_weights[34][33] = 16'sd6;
        fc1_weights[34][34] = 16'sd27;
        fc1_weights[34][35] = 16'sd20;
        fc1_weights[34][36] = 16'sd40;
        fc1_weights[34][37] = 16'sd60;
        fc1_weights[34][38] = 16'sd24;
        fc1_weights[34][39] = 16'sd-121;
        fc1_weights[34][40] = 16'sd26;
        fc1_weights[34][41] = 16'sd2;
        fc1_weights[34][42] = 16'sd-17;
        fc1_weights[34][43] = 16'sd20;
        fc1_weights[34][44] = 16'sd-28;
        fc1_weights[34][45] = 16'sd-26;
        fc1_weights[34][46] = 16'sd6;
        fc1_weights[34][47] = 16'sd-13;
        fc1_weights[34][48] = 16'sd1;
        fc1_weights[34][49] = 16'sd44;
        fc1_weights[34][50] = 16'sd-10;
        fc1_weights[34][51] = 16'sd6;
        fc1_weights[34][52] = 16'sd-53;
        fc1_weights[34][53] = 16'sd-43;
        fc1_weights[34][54] = 16'sd-2;
        fc1_weights[34][55] = 16'sd-36;
        fc1_weights[34][56] = 16'sd-42;
        fc1_weights[34][57] = 16'sd42;
        fc1_weights[34][58] = 16'sd23;
        fc1_weights[34][59] = 16'sd5;
        fc1_weights[34][60] = 16'sd37;
        fc1_weights[34][61] = 16'sd32;
        fc1_weights[34][62] = 16'sd16;
        fc1_weights[34][63] = 16'sd21;
        fc1_weights[34][64] = 16'sd-1;
        fc1_weights[34][65] = 16'sd18;
        fc1_weights[34][66] = 16'sd-30;
        fc1_weights[34][67] = 16'sd7;
        fc1_weights[34][68] = 16'sd-32;
        fc1_weights[34][69] = 16'sd-33;
        fc1_weights[34][70] = 16'sd-42;
        fc1_weights[34][71] = 16'sd-14;
        fc1_weights[34][72] = 16'sd7;
        fc1_weights[34][73] = 16'sd-34;
        fc1_weights[34][74] = 16'sd-12;
        fc1_weights[34][75] = 16'sd-21;
        fc1_weights[34][76] = 16'sd33;
        fc1_weights[34][77] = 16'sd-25;
        fc1_weights[34][78] = 16'sd35;
        fc1_weights[34][79] = 16'sd90;
        fc1_weights[34][80] = 16'sd-21;
        fc1_weights[34][81] = 16'sd3;
        fc1_weights[34][82] = 16'sd-40;
        fc1_weights[34][83] = 16'sd-9;
        fc1_weights[34][84] = 16'sd16;
        fc1_weights[34][85] = 16'sd-54;
        fc1_weights[34][86] = 16'sd-20;
        fc1_weights[34][87] = 16'sd0;
        fc1_weights[34][88] = 16'sd-66;
        fc1_weights[34][89] = 16'sd48;
        fc1_weights[34][90] = 16'sd-9;
        fc1_weights[34][91] = 16'sd-18;
        fc1_weights[34][92] = 16'sd-18;
        fc1_weights[34][93] = 16'sd-20;
        fc1_weights[34][94] = 16'sd-17;
        fc1_weights[34][95] = 16'sd0;
        fc1_weights[34][96] = 16'sd10;
        fc1_weights[34][97] = 16'sd-16;
        fc1_weights[34][98] = 16'sd-37;
        fc1_weights[34][99] = 16'sd-48;
        fc1_weights[34][100] = 16'sd16;
        fc1_weights[34][101] = 16'sd-13;
        fc1_weights[34][102] = 16'sd-38;
        fc1_weights[34][103] = 16'sd-47;
        fc1_weights[34][104] = 16'sd2;
        fc1_weights[34][105] = 16'sd-48;
        fc1_weights[34][106] = 16'sd-44;
        fc1_weights[34][107] = 16'sd-38;
        fc1_weights[34][108] = 16'sd1;
        fc1_weights[34][109] = 16'sd-14;
        fc1_weights[34][110] = 16'sd27;
        fc1_weights[34][111] = 16'sd-46;
        fc1_weights[34][112] = 16'sd-6;
        fc1_weights[34][113] = 16'sd53;
        fc1_weights[34][114] = 16'sd8;
        fc1_weights[34][115] = 16'sd38;
        fc1_weights[34][116] = 16'sd110;
        fc1_weights[34][117] = 16'sd57;
        fc1_weights[34][118] = 16'sd-8;
        fc1_weights[34][119] = 16'sd19;
        fc1_weights[34][120] = 16'sd28;
        fc1_weights[34][121] = 16'sd37;
        fc1_weights[34][122] = 16'sd16;
        fc1_weights[34][123] = 16'sd-17;
        fc1_weights[34][124] = 16'sd-35;
        fc1_weights[34][125] = 16'sd-7;
        fc1_weights[34][126] = 16'sd-37;
        fc1_weights[34][127] = 16'sd-38;
        fc1_weights[34][128] = 16'sd-25;
        fc1_weights[34][129] = 16'sd-48;
        fc1_weights[34][130] = 16'sd14;
        fc1_weights[34][131] = 16'sd-20;
        fc1_weights[34][132] = 16'sd-12;
        fc1_weights[34][133] = 16'sd-7;
        fc1_weights[34][134] = 16'sd4;
        fc1_weights[34][135] = 16'sd40;
        fc1_weights[34][136] = 16'sd15;
        fc1_weights[34][137] = 16'sd21;
        fc1_weights[34][138] = 16'sd-27;
        fc1_weights[34][139] = 16'sd15;
        fc1_weights[34][140] = 16'sd15;
        fc1_weights[34][141] = 16'sd-68;
        fc1_weights[34][142] = 16'sd2;
        fc1_weights[34][143] = 16'sd-21;
        fc1_weights[34][144] = 16'sd37;
        fc1_weights[34][145] = 16'sd1;
        fc1_weights[34][146] = 16'sd17;
        fc1_weights[34][147] = 16'sd36;
        fc1_weights[34][148] = 16'sd21;
        fc1_weights[34][149] = 16'sd12;
        fc1_weights[34][150] = 16'sd-77;
        fc1_weights[34][151] = 16'sd33;
        fc1_weights[34][152] = 16'sd1;
        fc1_weights[34][153] = 16'sd-25;
        fc1_weights[34][154] = 16'sd-5;
        fc1_weights[34][155] = 16'sd59;
        fc1_weights[34][156] = 16'sd20;
        fc1_weights[34][157] = 16'sd-7;
        fc1_weights[34][158] = 16'sd-22;
        fc1_weights[34][159] = 16'sd54;
        fc1_weights[34][160] = 16'sd-14;
        fc1_weights[34][161] = 16'sd3;
        fc1_weights[34][162] = 16'sd13;
        fc1_weights[34][163] = 16'sd-4;
        fc1_weights[34][164] = 16'sd-15;
        fc1_weights[34][165] = 16'sd24;
        fc1_weights[34][166] = 16'sd59;
        fc1_weights[34][167] = 16'sd19;
        fc1_weights[34][168] = 16'sd45;
        fc1_weights[34][169] = 16'sd-14;
        fc1_weights[34][170] = 16'sd10;
        fc1_weights[34][171] = 16'sd-3;
        fc1_weights[34][172] = 16'sd4;
        fc1_weights[34][173] = 16'sd-10;
        fc1_weights[34][174] = 16'sd11;
        fc1_weights[34][175] = 16'sd52;
        fc1_weights[34][176] = 16'sd26;
        fc1_weights[34][177] = 16'sd18;
        fc1_weights[34][178] = 16'sd21;
        fc1_weights[34][179] = 16'sd87;
        fc1_weights[34][180] = 16'sd63;
        fc1_weights[34][181] = 16'sd9;
        fc1_weights[34][182] = 16'sd14;
        fc1_weights[34][183] = 16'sd-3;
        fc1_weights[34][184] = 16'sd-7;
        fc1_weights[34][185] = 16'sd49;
        fc1_weights[34][186] = 16'sd-71;
        fc1_weights[34][187] = 16'sd5;
        fc1_weights[34][188] = 16'sd11;
        fc1_weights[34][189] = 16'sd-10;
        fc1_weights[34][190] = 16'sd105;
        fc1_weights[34][191] = 16'sd80;
        fc1_weights[34][192] = 16'sd-11;
        fc1_weights[34][193] = 16'sd25;
        fc1_weights[34][194] = 16'sd34;
        fc1_weights[34][195] = 16'sd-25;
        fc1_weights[34][196] = 16'sd-29;
        fc1_weights[34][197] = 16'sd35;
        fc1_weights[34][198] = 16'sd-7;
        fc1_weights[34][199] = 16'sd18;
        fc1_weights[34][200] = 16'sd1;
        fc1_weights[34][201] = 16'sd18;
        fc1_weights[34][202] = 16'sd-31;
        fc1_weights[34][203] = 16'sd57;
        fc1_weights[34][204] = 16'sd20;
        fc1_weights[34][205] = 16'sd68;
        fc1_weights[34][206] = 16'sd21;
        fc1_weights[34][207] = 16'sd14;
        fc1_weights[35][0] = 16'sd-32;
        fc1_weights[35][1] = 16'sd1;
        fc1_weights[35][2] = 16'sd-24;
        fc1_weights[35][3] = 16'sd-91;
        fc1_weights[35][4] = 16'sd-92;
        fc1_weights[35][5] = 16'sd-7;
        fc1_weights[35][6] = 16'sd-3;
        fc1_weights[35][7] = 16'sd-41;
        fc1_weights[35][8] = 16'sd-43;
        fc1_weights[35][9] = 16'sd23;
        fc1_weights[35][10] = 16'sd-17;
        fc1_weights[35][11] = 16'sd-125;
        fc1_weights[35][12] = 16'sd-178;
        fc1_weights[35][13] = 16'sd-43;
        fc1_weights[35][14] = 16'sd-34;
        fc1_weights[35][15] = 16'sd71;
        fc1_weights[35][16] = 16'sd-35;
        fc1_weights[35][17] = 16'sd-61;
        fc1_weights[35][18] = 16'sd-36;
        fc1_weights[35][19] = 16'sd4;
        fc1_weights[35][20] = 16'sd80;
        fc1_weights[35][21] = 16'sd14;
        fc1_weights[35][22] = 16'sd23;
        fc1_weights[35][23] = 16'sd-11;
        fc1_weights[35][24] = 16'sd42;
        fc1_weights[35][25] = 16'sd11;
        fc1_weights[35][26] = 16'sd-66;
        fc1_weights[35][27] = 16'sd34;
        fc1_weights[35][28] = 16'sd48;
        fc1_weights[35][29] = 16'sd-68;
        fc1_weights[35][30] = 16'sd-14;
        fc1_weights[35][31] = 16'sd-14;
        fc1_weights[35][32] = 16'sd5;
        fc1_weights[35][33] = 16'sd-59;
        fc1_weights[35][34] = 16'sd-54;
        fc1_weights[35][35] = 16'sd-60;
        fc1_weights[35][36] = 16'sd76;
        fc1_weights[35][37] = 16'sd-125;
        fc1_weights[35][38] = 16'sd-46;
        fc1_weights[35][39] = 16'sd-12;
        fc1_weights[35][40] = 16'sd110;
        fc1_weights[35][41] = 16'sd35;
        fc1_weights[35][42] = 16'sd-81;
        fc1_weights[35][43] = 16'sd18;
        fc1_weights[35][44] = 16'sd13;
        fc1_weights[35][45] = 16'sd-9;
        fc1_weights[35][46] = 16'sd-40;
        fc1_weights[35][47] = 16'sd-47;
        fc1_weights[35][48] = 16'sd18;
        fc1_weights[35][49] = 16'sd60;
        fc1_weights[35][50] = 16'sd32;
        fc1_weights[35][51] = 16'sd-89;
        fc1_weights[35][52] = 16'sd10;
        fc1_weights[35][53] = 16'sd58;
        fc1_weights[35][54] = 16'sd0;
        fc1_weights[35][55] = 16'sd31;
        fc1_weights[35][56] = 16'sd55;
        fc1_weights[35][57] = 16'sd42;
        fc1_weights[35][58] = 16'sd65;
        fc1_weights[35][59] = 16'sd9;
        fc1_weights[35][60] = 16'sd56;
        fc1_weights[35][61] = 16'sd52;
        fc1_weights[35][62] = 16'sd-30;
        fc1_weights[35][63] = 16'sd-3;
        fc1_weights[35][64] = 16'sd-15;
        fc1_weights[35][65] = 16'sd-99;
        fc1_weights[35][66] = 16'sd50;
        fc1_weights[35][67] = 16'sd25;
        fc1_weights[35][68] = 16'sd-20;
        fc1_weights[35][69] = 16'sd-57;
        fc1_weights[35][70] = 16'sd39;
        fc1_weights[35][71] = 16'sd40;
        fc1_weights[35][72] = 16'sd15;
        fc1_weights[35][73] = 16'sd-40;
        fc1_weights[35][74] = 16'sd-24;
        fc1_weights[35][75] = 16'sd20;
        fc1_weights[35][76] = 16'sd94;
        fc1_weights[35][77] = 16'sd16;
        fc1_weights[35][78] = 16'sd2;
        fc1_weights[35][79] = 16'sd97;
        fc1_weights[35][80] = 16'sd40;
        fc1_weights[35][81] = 16'sd47;
        fc1_weights[35][82] = 16'sd17;
        fc1_weights[35][83] = 16'sd-5;
        fc1_weights[35][84] = 16'sd-17;
        fc1_weights[35][85] = 16'sd-9;
        fc1_weights[35][86] = 16'sd55;
        fc1_weights[35][87] = 16'sd-11;
        fc1_weights[35][88] = 16'sd10;
        fc1_weights[35][89] = 16'sd-23;
        fc1_weights[35][90] = 16'sd78;
        fc1_weights[35][91] = 16'sd75;
        fc1_weights[35][92] = 16'sd1;
        fc1_weights[35][93] = 16'sd-24;
        fc1_weights[35][94] = 16'sd-9;
        fc1_weights[35][95] = 16'sd-30;
        fc1_weights[35][96] = 16'sd-4;
        fc1_weights[35][97] = 16'sd-46;
        fc1_weights[35][98] = 16'sd-37;
        fc1_weights[35][99] = 16'sd77;
        fc1_weights[35][100] = 16'sd16;
        fc1_weights[35][101] = 16'sd-13;
        fc1_weights[35][102] = 16'sd18;
        fc1_weights[35][103] = 16'sd-89;
        fc1_weights[35][104] = 16'sd-5;
        fc1_weights[35][105] = 16'sd-19;
        fc1_weights[35][106] = 16'sd-46;
        fc1_weights[35][107] = 16'sd44;
        fc1_weights[35][108] = 16'sd16;
        fc1_weights[35][109] = 16'sd21;
        fc1_weights[35][110] = 16'sd29;
        fc1_weights[35][111] = 16'sd-13;
        fc1_weights[35][112] = 16'sd69;
        fc1_weights[35][113] = 16'sd8;
        fc1_weights[35][114] = 16'sd-49;
        fc1_weights[35][115] = 16'sd-50;
        fc1_weights[35][116] = 16'sd-64;
        fc1_weights[35][117] = 16'sd50;
        fc1_weights[35][118] = 16'sd112;
        fc1_weights[35][119] = 16'sd37;
        fc1_weights[35][120] = 16'sd10;
        fc1_weights[35][121] = 16'sd-10;
        fc1_weights[35][122] = 16'sd30;
        fc1_weights[35][123] = 16'sd8;
        fc1_weights[35][124] = 16'sd-127;
        fc1_weights[35][125] = 16'sd28;
        fc1_weights[35][126] = 16'sd-52;
        fc1_weights[35][127] = 16'sd52;
        fc1_weights[35][128] = 16'sd-38;
        fc1_weights[35][129] = 16'sd-146;
        fc1_weights[35][130] = 16'sd-3;
        fc1_weights[35][131] = 16'sd11;
        fc1_weights[35][132] = 16'sd56;
        fc1_weights[35][133] = 16'sd48;
        fc1_weights[35][134] = 16'sd30;
        fc1_weights[35][135] = 16'sd65;
        fc1_weights[35][136] = 16'sd89;
        fc1_weights[35][137] = 16'sd94;
        fc1_weights[35][138] = 16'sd60;
        fc1_weights[35][139] = 16'sd-5;
        fc1_weights[35][140] = 16'sd-33;
        fc1_weights[35][141] = 16'sd-86;
        fc1_weights[35][142] = 16'sd7;
        fc1_weights[35][143] = 16'sd1;
        fc1_weights[35][144] = 16'sd7;
        fc1_weights[35][145] = 16'sd-37;
        fc1_weights[35][146] = 16'sd-47;
        fc1_weights[35][147] = 16'sd21;
        fc1_weights[35][148] = 16'sd17;
        fc1_weights[35][149] = 16'sd-33;
        fc1_weights[35][150] = 16'sd-18;
        fc1_weights[35][151] = 16'sd-9;
        fc1_weights[35][152] = 16'sd20;
        fc1_weights[35][153] = 16'sd83;
        fc1_weights[35][154] = 16'sd25;
        fc1_weights[35][155] = 16'sd25;
        fc1_weights[35][156] = 16'sd-22;
        fc1_weights[35][157] = 16'sd58;
        fc1_weights[35][158] = 16'sd27;
        fc1_weights[35][159] = 16'sd-87;
        fc1_weights[35][160] = 16'sd-87;
        fc1_weights[35][161] = 16'sd21;
        fc1_weights[35][162] = 16'sd12;
        fc1_weights[35][163] = 16'sd-5;
        fc1_weights[35][164] = 16'sd16;
        fc1_weights[35][165] = 16'sd-44;
        fc1_weights[35][166] = 16'sd-37;
        fc1_weights[35][167] = 16'sd26;
        fc1_weights[35][168] = 16'sd16;
        fc1_weights[35][169] = 16'sd37;
        fc1_weights[35][170] = 16'sd13;
        fc1_weights[35][171] = 16'sd32;
        fc1_weights[35][172] = 16'sd10;
        fc1_weights[35][173] = 16'sd1;
        fc1_weights[35][174] = 16'sd-40;
        fc1_weights[35][175] = 16'sd-14;
        fc1_weights[35][176] = 16'sd-68;
        fc1_weights[35][177] = 16'sd-43;
        fc1_weights[35][178] = 16'sd-67;
        fc1_weights[35][179] = 16'sd-64;
        fc1_weights[35][180] = 16'sd-46;
        fc1_weights[35][181] = 16'sd-2;
        fc1_weights[35][182] = 16'sd-51;
        fc1_weights[35][183] = 16'sd33;
        fc1_weights[35][184] = 16'sd10;
        fc1_weights[35][185] = 16'sd-2;
        fc1_weights[35][186] = 16'sd-38;
        fc1_weights[35][187] = 16'sd14;
        fc1_weights[35][188] = 16'sd-58;
        fc1_weights[35][189] = 16'sd-2;
        fc1_weights[35][190] = 16'sd-19;
        fc1_weights[35][191] = 16'sd42;
        fc1_weights[35][192] = 16'sd12;
        fc1_weights[35][193] = 16'sd48;
        fc1_weights[35][194] = 16'sd60;
        fc1_weights[35][195] = 16'sd36;
        fc1_weights[35][196] = 16'sd56;
        fc1_weights[35][197] = 16'sd106;
        fc1_weights[35][198] = 16'sd-38;
        fc1_weights[35][199] = 16'sd13;
        fc1_weights[35][200] = 16'sd42;
        fc1_weights[35][201] = 16'sd-7;
        fc1_weights[35][202] = 16'sd19;
        fc1_weights[35][203] = 16'sd8;
        fc1_weights[35][204] = 16'sd-7;
        fc1_weights[35][205] = 16'sd-33;
        fc1_weights[35][206] = 16'sd-28;
        fc1_weights[35][207] = 16'sd-68;
        fc1_weights[36][0] = 16'sd16;
        fc1_weights[36][1] = 16'sd10;
        fc1_weights[36][2] = 16'sd-4;
        fc1_weights[36][3] = 16'sd-12;
        fc1_weights[36][4] = 16'sd-26;
        fc1_weights[36][5] = 16'sd1;
        fc1_weights[36][6] = 16'sd51;
        fc1_weights[36][7] = 16'sd58;
        fc1_weights[36][8] = 16'sd8;
        fc1_weights[36][9] = 16'sd12;
        fc1_weights[36][10] = 16'sd-11;
        fc1_weights[36][11] = 16'sd-3;
        fc1_weights[36][12] = 16'sd10;
        fc1_weights[36][13] = 16'sd15;
        fc1_weights[36][14] = 16'sd8;
        fc1_weights[36][15] = 16'sd-40;
        fc1_weights[36][16] = 16'sd12;
        fc1_weights[36][17] = 16'sd11;
        fc1_weights[36][18] = 16'sd-13;
        fc1_weights[36][19] = 16'sd-20;
        fc1_weights[36][20] = 16'sd-5;
        fc1_weights[36][21] = 16'sd34;
        fc1_weights[36][22] = 16'sd14;
        fc1_weights[36][23] = 16'sd2;
        fc1_weights[36][24] = 16'sd33;
        fc1_weights[36][25] = 16'sd-8;
        fc1_weights[36][26] = 16'sd-9;
        fc1_weights[36][27] = 16'sd-6;
        fc1_weights[36][28] = 16'sd10;
        fc1_weights[36][29] = 16'sd-7;
        fc1_weights[36][30] = 16'sd0;
        fc1_weights[36][31] = 16'sd25;
        fc1_weights[36][32] = 16'sd10;
        fc1_weights[36][33] = 16'sd48;
        fc1_weights[36][34] = 16'sd94;
        fc1_weights[36][35] = 16'sd11;
        fc1_weights[36][36] = 16'sd-6;
        fc1_weights[36][37] = 16'sd40;
        fc1_weights[36][38] = 16'sd9;
        fc1_weights[36][39] = 16'sd-18;
        fc1_weights[36][40] = 16'sd23;
        fc1_weights[36][41] = 16'sd-15;
        fc1_weights[36][42] = 16'sd16;
        fc1_weights[36][43] = 16'sd-21;
        fc1_weights[36][44] = 16'sd-13;
        fc1_weights[36][45] = 16'sd27;
        fc1_weights[36][46] = 16'sd-9;
        fc1_weights[36][47] = 16'sd34;
        fc1_weights[36][48] = 16'sd5;
        fc1_weights[36][49] = 16'sd12;
        fc1_weights[36][50] = 16'sd32;
        fc1_weights[36][51] = 16'sd44;
        fc1_weights[36][52] = 16'sd11;
        fc1_weights[36][53] = 16'sd-36;
        fc1_weights[36][54] = 16'sd12;
        fc1_weights[36][55] = 16'sd25;
        fc1_weights[36][56] = 16'sd7;
        fc1_weights[36][57] = 16'sd10;
        fc1_weights[36][58] = 16'sd-18;
        fc1_weights[36][59] = 16'sd32;
        fc1_weights[36][60] = 16'sd24;
        fc1_weights[36][61] = 16'sd12;
        fc1_weights[36][62] = 16'sd3;
        fc1_weights[36][63] = 16'sd14;
        fc1_weights[36][64] = 16'sd36;
        fc1_weights[36][65] = 16'sd16;
        fc1_weights[36][66] = 16'sd47;
        fc1_weights[36][67] = 16'sd16;
        fc1_weights[36][68] = 16'sd-38;
        fc1_weights[36][69] = 16'sd14;
        fc1_weights[36][70] = 16'sd33;
        fc1_weights[36][71] = 16'sd37;
        fc1_weights[36][72] = 16'sd40;
        fc1_weights[36][73] = 16'sd46;
        fc1_weights[36][74] = 16'sd33;
        fc1_weights[36][75] = 16'sd33;
        fc1_weights[36][76] = 16'sd42;
        fc1_weights[36][77] = 16'sd83;
        fc1_weights[36][78] = 16'sd-9;
        fc1_weights[36][79] = 16'sd-8;
        fc1_weights[36][80] = 16'sd-29;
        fc1_weights[36][81] = 16'sd-16;
        fc1_weights[36][82] = 16'sd-55;
        fc1_weights[36][83] = 16'sd52;
        fc1_weights[36][84] = 16'sd10;
        fc1_weights[36][85] = 16'sd14;
        fc1_weights[36][86] = 16'sd17;
        fc1_weights[36][87] = 16'sd30;
        fc1_weights[36][88] = 16'sd33;
        fc1_weights[36][89] = 16'sd-4;
        fc1_weights[36][90] = 16'sd-36;
        fc1_weights[36][91] = 16'sd-8;
        fc1_weights[36][92] = 16'sd3;
        fc1_weights[36][93] = 16'sd6;
        fc1_weights[36][94] = 16'sd-25;
        fc1_weights[36][95] = 16'sd-16;
        fc1_weights[36][96] = 16'sd9;
        fc1_weights[36][97] = 16'sd39;
        fc1_weights[36][98] = 16'sd15;
        fc1_weights[36][99] = 16'sd24;
        fc1_weights[36][100] = 16'sd25;
        fc1_weights[36][101] = 16'sd32;
        fc1_weights[36][102] = 16'sd64;
        fc1_weights[36][103] = 16'sd70;
        fc1_weights[36][104] = 16'sd12;
        fc1_weights[36][105] = 16'sd1;
        fc1_weights[36][106] = 16'sd21;
        fc1_weights[36][107] = 16'sd25;
        fc1_weights[36][108] = 16'sd-13;
        fc1_weights[36][109] = 16'sd35;
        fc1_weights[36][110] = 16'sd-24;
        fc1_weights[36][111] = 16'sd-12;
        fc1_weights[36][112] = 16'sd-33;
        fc1_weights[36][113] = 16'sd-1;
        fc1_weights[36][114] = 16'sd40;
        fc1_weights[36][115] = 16'sd32;
        fc1_weights[36][116] = 16'sd-6;
        fc1_weights[36][117] = 16'sd-16;
        fc1_weights[36][118] = 16'sd-36;
        fc1_weights[36][119] = 16'sd-33;
        fc1_weights[36][120] = 16'sd-9;
        fc1_weights[36][121] = 16'sd3;
        fc1_weights[36][122] = 16'sd-6;
        fc1_weights[36][123] = 16'sd-15;
        fc1_weights[36][124] = 16'sd1;
        fc1_weights[36][125] = 16'sd14;
        fc1_weights[36][126] = 16'sd24;
        fc1_weights[36][127] = 16'sd-34;
        fc1_weights[36][128] = 16'sd-7;
        fc1_weights[36][129] = 16'sd47;
        fc1_weights[36][130] = 16'sd-5;
        fc1_weights[36][131] = 16'sd44;
        fc1_weights[36][132] = 16'sd41;
        fc1_weights[36][133] = 16'sd22;
        fc1_weights[36][134] = 16'sd-32;
        fc1_weights[36][135] = 16'sd31;
        fc1_weights[36][136] = 16'sd-1;
        fc1_weights[36][137] = 16'sd-2;
        fc1_weights[36][138] = 16'sd27;
        fc1_weights[36][139] = 16'sd-16;
        fc1_weights[36][140] = 16'sd20;
        fc1_weights[36][141] = 16'sd44;
        fc1_weights[36][142] = 16'sd-5;
        fc1_weights[36][143] = 16'sd-11;
        fc1_weights[36][144] = 16'sd23;
        fc1_weights[36][145] = 16'sd-10;
        fc1_weights[36][146] = 16'sd0;
        fc1_weights[36][147] = 16'sd-23;
        fc1_weights[36][148] = 16'sd23;
        fc1_weights[36][149] = 16'sd10;
        fc1_weights[36][150] = 16'sd35;
        fc1_weights[36][151] = 16'sd19;
        fc1_weights[36][152] = 16'sd-11;
        fc1_weights[36][153] = 16'sd-11;
        fc1_weights[36][154] = 16'sd-23;
        fc1_weights[36][155] = 16'sd1;
        fc1_weights[36][156] = 16'sd24;
        fc1_weights[36][157] = 16'sd-10;
        fc1_weights[36][158] = 16'sd41;
        fc1_weights[36][159] = 16'sd54;
        fc1_weights[36][160] = 16'sd14;
        fc1_weights[36][161] = 16'sd13;
        fc1_weights[36][162] = 16'sd9;
        fc1_weights[36][163] = 16'sd15;
        fc1_weights[36][164] = 16'sd-28;
        fc1_weights[36][165] = 16'sd21;
        fc1_weights[36][166] = 16'sd2;
        fc1_weights[36][167] = 16'sd9;
        fc1_weights[36][168] = 16'sd23;
        fc1_weights[36][169] = 16'sd2;
        fc1_weights[36][170] = 16'sd-13;
        fc1_weights[36][171] = 16'sd20;
        fc1_weights[36][172] = 16'sd-12;
        fc1_weights[36][173] = 16'sd1;
        fc1_weights[36][174] = 16'sd30;
        fc1_weights[36][175] = 16'sd7;
        fc1_weights[36][176] = 16'sd24;
        fc1_weights[36][177] = 16'sd18;
        fc1_weights[36][178] = 16'sd-3;
        fc1_weights[36][179] = 16'sd6;
        fc1_weights[36][180] = 16'sd49;
        fc1_weights[36][181] = 16'sd45;
        fc1_weights[36][182] = 16'sd37;
        fc1_weights[36][183] = 16'sd44;
        fc1_weights[36][184] = 16'sd13;
        fc1_weights[36][185] = 16'sd10;
        fc1_weights[36][186] = 16'sd-17;
        fc1_weights[36][187] = 16'sd-31;
        fc1_weights[36][188] = 16'sd-4;
        fc1_weights[36][189] = 16'sd-32;
        fc1_weights[36][190] = 16'sd-10;
        fc1_weights[36][191] = 16'sd8;
        fc1_weights[36][192] = 16'sd23;
        fc1_weights[36][193] = 16'sd-13;
        fc1_weights[36][194] = 16'sd-55;
        fc1_weights[36][195] = 16'sd-71;
        fc1_weights[36][196] = 16'sd-59;
        fc1_weights[36][197] = 16'sd-32;
        fc1_weights[36][198] = 16'sd-16;
        fc1_weights[36][199] = 16'sd-82;
        fc1_weights[36][200] = 16'sd-45;
        fc1_weights[36][201] = 16'sd-49;
        fc1_weights[36][202] = 16'sd-14;
        fc1_weights[36][203] = 16'sd-37;
        fc1_weights[36][204] = 16'sd-48;
        fc1_weights[36][205] = 16'sd-19;
        fc1_weights[36][206] = 16'sd1;
        fc1_weights[36][207] = 16'sd-8;
        fc1_weights[37][0] = 16'sd-10;
        fc1_weights[37][1] = 16'sd-8;
        fc1_weights[37][2] = 16'sd-1;
        fc1_weights[37][3] = 16'sd2;
        fc1_weights[37][4] = 16'sd9;
        fc1_weights[37][5] = 16'sd-10;
        fc1_weights[37][6] = 16'sd-6;
        fc1_weights[37][7] = 16'sd-5;
        fc1_weights[37][8] = 16'sd-20;
        fc1_weights[37][9] = 16'sd5;
        fc1_weights[37][10] = 16'sd8;
        fc1_weights[37][11] = 16'sd14;
        fc1_weights[37][12] = 16'sd29;
        fc1_weights[37][13] = 16'sd21;
        fc1_weights[37][14] = 16'sd-8;
        fc1_weights[37][15] = 16'sd-24;
        fc1_weights[37][16] = 16'sd24;
        fc1_weights[37][17] = 16'sd34;
        fc1_weights[37][18] = 16'sd63;
        fc1_weights[37][19] = 16'sd65;
        fc1_weights[37][20] = 16'sd54;
        fc1_weights[37][21] = 16'sd48;
        fc1_weights[37][22] = 16'sd9;
        fc1_weights[37][23] = 16'sd-10;
        fc1_weights[37][24] = 16'sd13;
        fc1_weights[37][25] = 16'sd9;
        fc1_weights[37][26] = 16'sd-32;
        fc1_weights[37][27] = 16'sd-13;
        fc1_weights[37][28] = 16'sd-43;
        fc1_weights[37][29] = 16'sd-18;
        fc1_weights[37][30] = 16'sd18;
        fc1_weights[37][31] = 16'sd-9;
        fc1_weights[37][32] = 16'sd-32;
        fc1_weights[37][33] = 16'sd49;
        fc1_weights[37][34] = 16'sd4;
        fc1_weights[37][35] = 16'sd-6;
        fc1_weights[37][36] = 16'sd-34;
        fc1_weights[37][37] = 16'sd18;
        fc1_weights[37][38] = 16'sd41;
        fc1_weights[37][39] = 16'sd51;
        fc1_weights[37][40] = 16'sd3;
        fc1_weights[37][41] = 16'sd21;
        fc1_weights[37][42] = 16'sd71;
        fc1_weights[37][43] = 16'sd40;
        fc1_weights[37][44] = 16'sd48;
        fc1_weights[37][45] = 16'sd21;
        fc1_weights[37][46] = 16'sd26;
        fc1_weights[37][47] = 16'sd7;
        fc1_weights[37][48] = 16'sd11;
        fc1_weights[37][49] = 16'sd16;
        fc1_weights[37][50] = 16'sd2;
        fc1_weights[37][51] = 16'sd31;
        fc1_weights[37][52] = 16'sd-18;
        fc1_weights[37][53] = 16'sd-25;
        fc1_weights[37][54] = 16'sd4;
        fc1_weights[37][55] = 16'sd-68;
        fc1_weights[37][56] = 16'sd-42;
        fc1_weights[37][57] = 16'sd-13;
        fc1_weights[37][58] = 16'sd6;
        fc1_weights[37][59] = 16'sd-1;
        fc1_weights[37][60] = 16'sd-8;
        fc1_weights[37][61] = 16'sd3;
        fc1_weights[37][62] = 16'sd80;
        fc1_weights[37][63] = 16'sd6;
        fc1_weights[37][64] = 16'sd15;
        fc1_weights[37][65] = 16'sd33;
        fc1_weights[37][66] = 16'sd26;
        fc1_weights[37][67] = 16'sd33;
        fc1_weights[37][68] = 16'sd38;
        fc1_weights[37][69] = 16'sd-8;
        fc1_weights[37][70] = 16'sd-23;
        fc1_weights[37][71] = 16'sd28;
        fc1_weights[37][72] = 16'sd10;
        fc1_weights[37][73] = 16'sd11;
        fc1_weights[37][74] = 16'sd3;
        fc1_weights[37][75] = 16'sd13;
        fc1_weights[37][76] = 16'sd3;
        fc1_weights[37][77] = 16'sd41;
        fc1_weights[37][78] = 16'sd60;
        fc1_weights[37][79] = 16'sd2;
        fc1_weights[37][80] = 16'sd35;
        fc1_weights[37][81] = 16'sd-7;
        fc1_weights[37][82] = 16'sd29;
        fc1_weights[37][83] = 16'sd-2;
        fc1_weights[37][84] = 16'sd5;
        fc1_weights[37][85] = 16'sd-9;
        fc1_weights[37][86] = 16'sd10;
        fc1_weights[37][87] = 16'sd-36;
        fc1_weights[37][88] = 16'sd-12;
        fc1_weights[37][89] = 16'sd-17;
        fc1_weights[37][90] = 16'sd-5;
        fc1_weights[37][91] = 16'sd13;
        fc1_weights[37][92] = 16'sd-67;
        fc1_weights[37][93] = 16'sd-67;
        fc1_weights[37][94] = 16'sd36;
        fc1_weights[37][95] = 16'sd-22;
        fc1_weights[37][96] = 16'sd-25;
        fc1_weights[37][97] = 16'sd28;
        fc1_weights[37][98] = 16'sd-32;
        fc1_weights[37][99] = 16'sd24;
        fc1_weights[37][100] = 16'sd-5;
        fc1_weights[37][101] = 16'sd13;
        fc1_weights[37][102] = 16'sd1;
        fc1_weights[37][103] = 16'sd8;
        fc1_weights[37][104] = 16'sd-16;
        fc1_weights[37][105] = 16'sd32;
        fc1_weights[37][106] = 16'sd-43;
        fc1_weights[37][107] = 16'sd-49;
        fc1_weights[37][108] = 16'sd24;
        fc1_weights[37][109] = 16'sd1;
        fc1_weights[37][110] = 16'sd-7;
        fc1_weights[37][111] = 16'sd-31;
        fc1_weights[37][112] = 16'sd-11;
        fc1_weights[37][113] = 16'sd6;
        fc1_weights[37][114] = 16'sd29;
        fc1_weights[37][115] = 16'sd24;
        fc1_weights[37][116] = 16'sd-10;
        fc1_weights[37][117] = 16'sd-27;
        fc1_weights[37][118] = 16'sd-19;
        fc1_weights[37][119] = 16'sd-18;
        fc1_weights[37][120] = 16'sd0;
        fc1_weights[37][121] = 16'sd-43;
        fc1_weights[37][122] = 16'sd-35;
        fc1_weights[37][123] = 16'sd-16;
        fc1_weights[37][124] = 16'sd-3;
        fc1_weights[37][125] = 16'sd5;
        fc1_weights[37][126] = 16'sd21;
        fc1_weights[37][127] = 16'sd11;
        fc1_weights[37][128] = 16'sd-12;
        fc1_weights[37][129] = 16'sd-8;
        fc1_weights[37][130] = 16'sd19;
        fc1_weights[37][131] = 16'sd-26;
        fc1_weights[37][132] = 16'sd-10;
        fc1_weights[37][133] = 16'sd-14;
        fc1_weights[37][134] = 16'sd19;
        fc1_weights[37][135] = 16'sd-4;
        fc1_weights[37][136] = 16'sd-7;
        fc1_weights[37][137] = 16'sd29;
        fc1_weights[37][138] = 16'sd21;
        fc1_weights[37][139] = 16'sd30;
        fc1_weights[37][140] = 16'sd25;
        fc1_weights[37][141] = 16'sd0;
        fc1_weights[37][142] = 16'sd-62;
        fc1_weights[37][143] = 16'sd-41;
        fc1_weights[37][144] = 16'sd-33;
        fc1_weights[37][145] = 16'sd-39;
        fc1_weights[37][146] = 16'sd-28;
        fc1_weights[37][147] = 16'sd-36;
        fc1_weights[37][148] = 16'sd-19;
        fc1_weights[37][149] = 16'sd2;
        fc1_weights[37][150] = 16'sd-24;
        fc1_weights[37][151] = 16'sd-32;
        fc1_weights[37][152] = 16'sd-26;
        fc1_weights[37][153] = 16'sd-47;
        fc1_weights[37][154] = 16'sd-42;
        fc1_weights[37][155] = 16'sd-3;
        fc1_weights[37][156] = 16'sd37;
        fc1_weights[37][157] = 16'sd11;
        fc1_weights[37][158] = 16'sd-4;
        fc1_weights[37][159] = 16'sd30;
        fc1_weights[37][160] = 16'sd21;
        fc1_weights[37][161] = 16'sd24;
        fc1_weights[37][162] = 16'sd15;
        fc1_weights[37][163] = 16'sd18;
        fc1_weights[37][164] = 16'sd37;
        fc1_weights[37][165] = 16'sd37;
        fc1_weights[37][166] = 16'sd33;
        fc1_weights[37][167] = 16'sd9;
        fc1_weights[37][168] = 16'sd23;
        fc1_weights[37][169] = 16'sd13;
        fc1_weights[37][170] = 16'sd9;
        fc1_weights[37][171] = 16'sd62;
        fc1_weights[37][172] = 16'sd8;
        fc1_weights[37][173] = 16'sd34;
        fc1_weights[37][174] = 16'sd21;
        fc1_weights[37][175] = 16'sd14;
        fc1_weights[37][176] = 16'sd-3;
        fc1_weights[37][177] = 16'sd8;
        fc1_weights[37][178] = 16'sd25;
        fc1_weights[37][179] = 16'sd-15;
        fc1_weights[37][180] = 16'sd-27;
        fc1_weights[37][181] = 16'sd-46;
        fc1_weights[37][182] = 16'sd60;
        fc1_weights[37][183] = 16'sd33;
        fc1_weights[37][184] = 16'sd48;
        fc1_weights[37][185] = 16'sd-1;
        fc1_weights[37][186] = 16'sd23;
        fc1_weights[37][187] = 16'sd35;
        fc1_weights[37][188] = 16'sd38;
        fc1_weights[37][189] = 16'sd28;
        fc1_weights[37][190] = 16'sd20;
        fc1_weights[37][191] = 16'sd24;
        fc1_weights[37][192] = 16'sd13;
        fc1_weights[37][193] = 16'sd26;
        fc1_weights[37][194] = 16'sd-3;
        fc1_weights[37][195] = 16'sd6;
        fc1_weights[37][196] = 16'sd-6;
        fc1_weights[37][197] = 16'sd5;
        fc1_weights[37][198] = 16'sd31;
        fc1_weights[37][199] = 16'sd-9;
        fc1_weights[37][200] = 16'sd-13;
        fc1_weights[37][201] = 16'sd10;
        fc1_weights[37][202] = 16'sd7;
        fc1_weights[37][203] = 16'sd-27;
        fc1_weights[37][204] = 16'sd0;
        fc1_weights[37][205] = 16'sd-31;
        fc1_weights[37][206] = 16'sd-35;
        fc1_weights[37][207] = 16'sd-41;
        fc1_weights[38][0] = 16'sd-42;
        fc1_weights[38][1] = 16'sd-8;
        fc1_weights[38][2] = 16'sd-21;
        fc1_weights[38][3] = 16'sd-69;
        fc1_weights[38][4] = 16'sd-75;
        fc1_weights[38][5] = 16'sd21;
        fc1_weights[38][6] = 16'sd-56;
        fc1_weights[38][7] = 16'sd-62;
        fc1_weights[38][8] = 16'sd-24;
        fc1_weights[38][9] = 16'sd1;
        fc1_weights[38][10] = 16'sd53;
        fc1_weights[38][11] = 16'sd44;
        fc1_weights[38][12] = 16'sd29;
        fc1_weights[38][13] = 16'sd29;
        fc1_weights[38][14] = 16'sd16;
        fc1_weights[38][15] = 16'sd2;
        fc1_weights[38][16] = 16'sd7;
        fc1_weights[38][17] = 16'sd43;
        fc1_weights[38][18] = 16'sd-10;
        fc1_weights[38][19] = 16'sd-52;
        fc1_weights[38][20] = 16'sd-81;
        fc1_weights[38][21] = 16'sd-27;
        fc1_weights[38][22] = 16'sd-90;
        fc1_weights[38][23] = 16'sd-2;
        fc1_weights[38][24] = 16'sd-46;
        fc1_weights[38][25] = 16'sd-1;
        fc1_weights[38][26] = 16'sd-20;
        fc1_weights[38][27] = 16'sd-22;
        fc1_weights[38][28] = 16'sd34;
        fc1_weights[38][29] = 16'sd1;
        fc1_weights[38][30] = 16'sd-32;
        fc1_weights[38][31] = 16'sd26;
        fc1_weights[38][32] = 16'sd-21;
        fc1_weights[38][33] = 16'sd-135;
        fc1_weights[38][34] = 16'sd-27;
        fc1_weights[38][35] = 16'sd-36;
        fc1_weights[38][36] = 16'sd-12;
        fc1_weights[38][37] = 16'sd22;
        fc1_weights[38][38] = 16'sd-31;
        fc1_weights[38][39] = 16'sd27;
        fc1_weights[38][40] = 16'sd-22;
        fc1_weights[38][41] = 16'sd-63;
        fc1_weights[38][42] = 16'sd-23;
        fc1_weights[38][43] = 16'sd-54;
        fc1_weights[38][44] = 16'sd-23;
        fc1_weights[38][45] = 16'sd-37;
        fc1_weights[38][46] = 16'sd-94;
        fc1_weights[38][47] = 16'sd-25;
        fc1_weights[38][48] = 16'sd-66;
        fc1_weights[38][49] = 16'sd-10;
        fc1_weights[38][50] = 16'sd39;
        fc1_weights[38][51] = 16'sd4;
        fc1_weights[38][52] = 16'sd40;
        fc1_weights[38][53] = 16'sd54;
        fc1_weights[38][54] = 16'sd31;
        fc1_weights[38][55] = 16'sd32;
        fc1_weights[38][56] = 16'sd16;
        fc1_weights[38][57] = 16'sd35;
        fc1_weights[38][58] = 16'sd28;
        fc1_weights[38][59] = 16'sd-26;
        fc1_weights[38][60] = 16'sd13;
        fc1_weights[38][61] = 16'sd-22;
        fc1_weights[38][62] = 16'sd10;
        fc1_weights[38][63] = 16'sd-10;
        fc1_weights[38][64] = 16'sd-19;
        fc1_weights[38][65] = 16'sd24;
        fc1_weights[38][66] = 16'sd13;
        fc1_weights[38][67] = 16'sd-35;
        fc1_weights[38][68] = 16'sd-67;
        fc1_weights[38][69] = 16'sd6;
        fc1_weights[38][70] = 16'sd71;
        fc1_weights[38][71] = 16'sd33;
        fc1_weights[38][72] = 16'sd-39;
        fc1_weights[38][73] = 16'sd3;
        fc1_weights[38][74] = 16'sd29;
        fc1_weights[38][75] = 16'sd-6;
        fc1_weights[38][76] = 16'sd-16;
        fc1_weights[38][77] = 16'sd18;
        fc1_weights[38][78] = 16'sd-42;
        fc1_weights[38][79] = 16'sd-32;
        fc1_weights[38][80] = 16'sd-6;
        fc1_weights[38][81] = 16'sd26;
        fc1_weights[38][82] = 16'sd-30;
        fc1_weights[38][83] = 16'sd46;
        fc1_weights[38][84] = 16'sd12;
        fc1_weights[38][85] = 16'sd19;
        fc1_weights[38][86] = 16'sd59;
        fc1_weights[38][87] = 16'sd74;
        fc1_weights[38][88] = 16'sd101;
        fc1_weights[38][89] = 16'sd-41;
        fc1_weights[38][90] = 16'sd-2;
        fc1_weights[38][91] = 16'sd-16;
        fc1_weights[38][92] = 16'sd36;
        fc1_weights[38][93] = 16'sd-41;
        fc1_weights[38][94] = 16'sd-50;
        fc1_weights[38][95] = 16'sd5;
        fc1_weights[38][96] = 16'sd-4;
        fc1_weights[38][97] = 16'sd17;
        fc1_weights[38][98] = 16'sd40;
        fc1_weights[38][99] = 16'sd-28;
        fc1_weights[38][100] = 16'sd-38;
        fc1_weights[38][101] = 16'sd-23;
        fc1_weights[38][102] = 16'sd-26;
        fc1_weights[38][103] = 16'sd20;
        fc1_weights[38][104] = 16'sd72;
        fc1_weights[38][105] = 16'sd11;
        fc1_weights[38][106] = 16'sd82;
        fc1_weights[38][107] = 16'sd61;
        fc1_weights[38][108] = 16'sd36;
        fc1_weights[38][109] = 16'sd-6;
        fc1_weights[38][110] = 16'sd-14;
        fc1_weights[38][111] = 16'sd43;
        fc1_weights[38][112] = 16'sd49;
        fc1_weights[38][113] = 16'sd17;
        fc1_weights[38][114] = 16'sd22;
        fc1_weights[38][115] = 16'sd77;
        fc1_weights[38][116] = 16'sd7;
        fc1_weights[38][117] = 16'sd6;
        fc1_weights[38][118] = 16'sd77;
        fc1_weights[38][119] = 16'sd-23;
        fc1_weights[38][120] = 16'sd37;
        fc1_weights[38][121] = 16'sd-4;
        fc1_weights[38][122] = 16'sd-10;
        fc1_weights[38][123] = 16'sd-11;
        fc1_weights[38][124] = 16'sd-68;
        fc1_weights[38][125] = 16'sd-78;
        fc1_weights[38][126] = 16'sd-13;
        fc1_weights[38][127] = 16'sd-30;
        fc1_weights[38][128] = 16'sd-15;
        fc1_weights[38][129] = 16'sd42;
        fc1_weights[38][130] = 16'sd-35;
        fc1_weights[38][131] = 16'sd-41;
        fc1_weights[38][132] = 16'sd-3;
        fc1_weights[38][133] = 16'sd-7;
        fc1_weights[38][134] = 16'sd-31;
        fc1_weights[38][135] = 16'sd-23;
        fc1_weights[38][136] = 16'sd-31;
        fc1_weights[38][137] = 16'sd-12;
        fc1_weights[38][138] = 16'sd25;
        fc1_weights[38][139] = 16'sd-73;
        fc1_weights[38][140] = 16'sd-55;
        fc1_weights[38][141] = 16'sd86;
        fc1_weights[38][142] = 16'sd6;
        fc1_weights[38][143] = 16'sd4;
        fc1_weights[38][144] = 16'sd22;
        fc1_weights[38][145] = 16'sd31;
        fc1_weights[38][146] = 16'sd28;
        fc1_weights[38][147] = 16'sd3;
        fc1_weights[38][148] = 16'sd-65;
        fc1_weights[38][149] = 16'sd-67;
        fc1_weights[38][150] = 16'sd-15;
        fc1_weights[38][151] = 16'sd-22;
        fc1_weights[38][152] = 16'sd-18;
        fc1_weights[38][153] = 16'sd-24;
        fc1_weights[38][154] = 16'sd-57;
        fc1_weights[38][155] = 16'sd7;
        fc1_weights[38][156] = 16'sd-54;
        fc1_weights[38][157] = 16'sd-35;
        fc1_weights[38][158] = 16'sd-10;
        fc1_weights[38][159] = 16'sd21;
        fc1_weights[38][160] = 16'sd20;
        fc1_weights[38][161] = 16'sd38;
        fc1_weights[38][162] = 16'sd72;
        fc1_weights[38][163] = 16'sd19;
        fc1_weights[38][164] = 16'sd-62;
        fc1_weights[38][165] = 16'sd-62;
        fc1_weights[38][166] = 16'sd-102;
        fc1_weights[38][167] = 16'sd-70;
        fc1_weights[38][168] = 16'sd-59;
        fc1_weights[38][169] = 16'sd-25;
        fc1_weights[38][170] = 16'sd42;
        fc1_weights[38][171] = 16'sd-40;
        fc1_weights[38][172] = 16'sd30;
        fc1_weights[38][173] = 16'sd-32;
        fc1_weights[38][174] = 16'sd7;
        fc1_weights[38][175] = 16'sd-38;
        fc1_weights[38][176] = 16'sd-39;
        fc1_weights[38][177] = 16'sd1;
        fc1_weights[38][178] = 16'sd28;
        fc1_weights[38][179] = 16'sd-38;
        fc1_weights[38][180] = 16'sd-5;
        fc1_weights[38][181] = 16'sd26;
        fc1_weights[38][182] = 16'sd-10;
        fc1_weights[38][183] = 16'sd-10;
        fc1_weights[38][184] = 16'sd-1;
        fc1_weights[38][185] = 16'sd-39;
        fc1_weights[38][186] = 16'sd52;
        fc1_weights[38][187] = 16'sd-45;
        fc1_weights[38][188] = 16'sd-28;
        fc1_weights[38][189] = 16'sd12;
        fc1_weights[38][190] = 16'sd23;
        fc1_weights[38][191] = 16'sd8;
        fc1_weights[38][192] = 16'sd50;
        fc1_weights[38][193] = 16'sd17;
        fc1_weights[38][194] = 16'sd8;
        fc1_weights[38][195] = 16'sd42;
        fc1_weights[38][196] = 16'sd55;
        fc1_weights[38][197] = 16'sd43;
        fc1_weights[38][198] = 16'sd-5;
        fc1_weights[38][199] = 16'sd49;
        fc1_weights[38][200] = 16'sd49;
        fc1_weights[38][201] = 16'sd14;
        fc1_weights[38][202] = 16'sd-32;
        fc1_weights[38][203] = 16'sd14;
        fc1_weights[38][204] = 16'sd-4;
        fc1_weights[38][205] = 16'sd-40;
        fc1_weights[38][206] = 16'sd21;
        fc1_weights[38][207] = 16'sd102;
        fc1_weights[39][0] = 16'sd63;
        fc1_weights[39][1] = 16'sd-27;
        fc1_weights[39][2] = 16'sd-20;
        fc1_weights[39][3] = 16'sd-25;
        fc1_weights[39][4] = 16'sd-30;
        fc1_weights[39][5] = 16'sd-61;
        fc1_weights[39][6] = 16'sd-20;
        fc1_weights[39][7] = 16'sd-16;
        fc1_weights[39][8] = 16'sd0;
        fc1_weights[39][9] = 16'sd-16;
        fc1_weights[39][10] = 16'sd-90;
        fc1_weights[39][11] = 16'sd59;
        fc1_weights[39][12] = 16'sd126;
        fc1_weights[39][13] = 16'sd46;
        fc1_weights[39][14] = 16'sd62;
        fc1_weights[39][15] = 16'sd-3;
        fc1_weights[39][16] = 16'sd3;
        fc1_weights[39][17] = 16'sd31;
        fc1_weights[39][18] = 16'sd11;
        fc1_weights[39][19] = 16'sd50;
        fc1_weights[39][20] = 16'sd13;
        fc1_weights[39][21] = 16'sd-6;
        fc1_weights[39][22] = 16'sd-69;
        fc1_weights[39][23] = 16'sd14;
        fc1_weights[39][24] = 16'sd-44;
        fc1_weights[39][25] = 16'sd-60;
        fc1_weights[39][26] = 16'sd56;
        fc1_weights[39][27] = 16'sd-11;
        fc1_weights[39][28] = 16'sd-31;
        fc1_weights[39][29] = 16'sd-41;
        fc1_weights[39][30] = 16'sd-19;
        fc1_weights[39][31] = 16'sd-40;
        fc1_weights[39][32] = 16'sd-1;
        fc1_weights[39][33] = 16'sd29;
        fc1_weights[39][34] = 16'sd38;
        fc1_weights[39][35] = 16'sd-6;
        fc1_weights[39][36] = 16'sd-65;
        fc1_weights[39][37] = 16'sd-6;
        fc1_weights[39][38] = 16'sd31;
        fc1_weights[39][39] = 16'sd-15;
        fc1_weights[39][40] = 16'sd-2;
        fc1_weights[39][41] = 16'sd8;
        fc1_weights[39][42] = 16'sd28;
        fc1_weights[39][43] = 16'sd-14;
        fc1_weights[39][44] = 16'sd-25;
        fc1_weights[39][45] = 16'sd37;
        fc1_weights[39][46] = 16'sd82;
        fc1_weights[39][47] = 16'sd12;
        fc1_weights[39][48] = 16'sd-3;
        fc1_weights[39][49] = 16'sd-19;
        fc1_weights[39][50] = 16'sd-16;
        fc1_weights[39][51] = 16'sd-12;
        fc1_weights[39][52] = 16'sd37;
        fc1_weights[39][53] = 16'sd-20;
        fc1_weights[39][54] = 16'sd-28;
        fc1_weights[39][55] = 16'sd0;
        fc1_weights[39][56] = 16'sd10;
        fc1_weights[39][57] = 16'sd-2;
        fc1_weights[39][58] = 16'sd36;
        fc1_weights[39][59] = 16'sd55;
        fc1_weights[39][60] = 16'sd17;
        fc1_weights[39][61] = 16'sd18;
        fc1_weights[39][62] = 16'sd70;
        fc1_weights[39][63] = 16'sd-22;
        fc1_weights[39][64] = 16'sd-64;
        fc1_weights[39][65] = 16'sd-7;
        fc1_weights[39][66] = 16'sd-24;
        fc1_weights[39][67] = 16'sd-37;
        fc1_weights[39][68] = 16'sd-80;
        fc1_weights[39][69] = 16'sd12;
        fc1_weights[39][70] = 16'sd30;
        fc1_weights[39][71] = 16'sd52;
        fc1_weights[39][72] = 16'sd20;
        fc1_weights[39][73] = 16'sd2;
        fc1_weights[39][74] = 16'sd-19;
        fc1_weights[39][75] = 16'sd1;
        fc1_weights[39][76] = 16'sd-9;
        fc1_weights[39][77] = 16'sd11;
        fc1_weights[39][78] = 16'sd-45;
        fc1_weights[39][79] = 16'sd-83;
        fc1_weights[39][80] = 16'sd-62;
        fc1_weights[39][81] = 16'sd-28;
        fc1_weights[39][82] = 16'sd-39;
        fc1_weights[39][83] = 16'sd-18;
        fc1_weights[39][84] = 16'sd43;
        fc1_weights[39][85] = 16'sd20;
        fc1_weights[39][86] = 16'sd-3;
        fc1_weights[39][87] = 16'sd-33;
        fc1_weights[39][88] = 16'sd3;
        fc1_weights[39][89] = 16'sd50;
        fc1_weights[39][90] = 16'sd-9;
        fc1_weights[39][91] = 16'sd-52;
        fc1_weights[39][92] = 16'sd13;
        fc1_weights[39][93] = 16'sd-38;
        fc1_weights[39][94] = 16'sd-39;
        fc1_weights[39][95] = 16'sd-54;
        fc1_weights[39][96] = 16'sd54;
        fc1_weights[39][97] = 16'sd14;
        fc1_weights[39][98] = 16'sd23;
        fc1_weights[39][99] = 16'sd-11;
        fc1_weights[39][100] = 16'sd12;
        fc1_weights[39][101] = 16'sd58;
        fc1_weights[39][102] = 16'sd25;
        fc1_weights[39][103] = 16'sd37;
        fc1_weights[39][104] = 16'sd-3;
        fc1_weights[39][105] = 16'sd27;
        fc1_weights[39][106] = 16'sd25;
        fc1_weights[39][107] = 16'sd-13;
        fc1_weights[39][108] = 16'sd-20;
        fc1_weights[39][109] = 16'sd8;
        fc1_weights[39][110] = 16'sd3;
        fc1_weights[39][111] = 16'sd-29;
        fc1_weights[39][112] = 16'sd-36;
        fc1_weights[39][113] = 16'sd50;
        fc1_weights[39][114] = 16'sd12;
        fc1_weights[39][115] = 16'sd88;
        fc1_weights[39][116] = 16'sd6;
        fc1_weights[39][117] = 16'sd-38;
        fc1_weights[39][118] = 16'sd-59;
        fc1_weights[39][119] = 16'sd-29;
        fc1_weights[39][120] = 16'sd-56;
        fc1_weights[39][121] = 16'sd-63;
        fc1_weights[39][122] = 16'sd-55;
        fc1_weights[39][123] = 16'sd-74;
        fc1_weights[39][124] = 16'sd49;
        fc1_weights[39][125] = 16'sd-44;
        fc1_weights[39][126] = 16'sd46;
        fc1_weights[39][127] = 16'sd-5;
        fc1_weights[39][128] = 16'sd6;
        fc1_weights[39][129] = 16'sd26;
        fc1_weights[39][130] = 16'sd38;
        fc1_weights[39][131] = 16'sd-8;
        fc1_weights[39][132] = 16'sd-5;
        fc1_weights[39][133] = 16'sd35;
        fc1_weights[39][134] = 16'sd-19;
        fc1_weights[39][135] = 16'sd-16;
        fc1_weights[39][136] = 16'sd14;
        fc1_weights[39][137] = 16'sd8;
        fc1_weights[39][138] = 16'sd36;
        fc1_weights[39][139] = 16'sd-15;
        fc1_weights[39][140] = 16'sd-5;
        fc1_weights[39][141] = 16'sd81;
        fc1_weights[39][142] = 16'sd16;
        fc1_weights[39][143] = 16'sd22;
        fc1_weights[39][144] = 16'sd35;
        fc1_weights[39][145] = 16'sd44;
        fc1_weights[39][146] = 16'sd19;
        fc1_weights[39][147] = 16'sd-3;
        fc1_weights[39][148] = 16'sd19;
        fc1_weights[39][149] = 16'sd29;
        fc1_weights[39][150] = 16'sd37;
        fc1_weights[39][151] = 16'sd-52;
        fc1_weights[39][152] = 16'sd-14;
        fc1_weights[39][153] = 16'sd-9;
        fc1_weights[39][154] = 16'sd6;
        fc1_weights[39][155] = 16'sd13;
        fc1_weights[39][156] = 16'sd-55;
        fc1_weights[39][157] = 16'sd-39;
        fc1_weights[39][158] = 16'sd16;
        fc1_weights[39][159] = 16'sd-6;
        fc1_weights[39][160] = 16'sd20;
        fc1_weights[39][161] = 16'sd28;
        fc1_weights[39][162] = 16'sd9;
        fc1_weights[39][163] = 16'sd-28;
        fc1_weights[39][164] = 16'sd14;
        fc1_weights[39][165] = 16'sd21;
        fc1_weights[39][166] = 16'sd-12;
        fc1_weights[39][167] = 16'sd26;
        fc1_weights[39][168] = 16'sd74;
        fc1_weights[39][169] = 16'sd86;
        fc1_weights[39][170] = 16'sd71;
        fc1_weights[39][171] = 16'sd104;
        fc1_weights[39][172] = 16'sd11;
        fc1_weights[39][173] = 16'sd-16;
        fc1_weights[39][174] = 16'sd-19;
        fc1_weights[39][175] = 16'sd-13;
        fc1_weights[39][176] = 16'sd-104;
        fc1_weights[39][177] = 16'sd-108;
        fc1_weights[39][178] = 16'sd-46;
        fc1_weights[39][179] = 16'sd-97;
        fc1_weights[39][180] = 16'sd-47;
        fc1_weights[39][181] = 16'sd-23;
        fc1_weights[39][182] = 16'sd-3;
        fc1_weights[39][183] = 16'sd-31;
        fc1_weights[39][184] = 16'sd-36;
        fc1_weights[39][185] = 16'sd-18;
        fc1_weights[39][186] = 16'sd28;
        fc1_weights[39][187] = 16'sd-22;
        fc1_weights[39][188] = 16'sd26;
        fc1_weights[39][189] = 16'sd60;
        fc1_weights[39][190] = 16'sd62;
        fc1_weights[39][191] = 16'sd-14;
        fc1_weights[39][192] = 16'sd2;
        fc1_weights[39][193] = 16'sd20;
        fc1_weights[39][194] = 16'sd30;
        fc1_weights[39][195] = 16'sd37;
        fc1_weights[39][196] = 16'sd33;
        fc1_weights[39][197] = 16'sd-6;
        fc1_weights[39][198] = 16'sd40;
        fc1_weights[39][199] = 16'sd10;
        fc1_weights[39][200] = 16'sd-31;
        fc1_weights[39][201] = 16'sd2;
        fc1_weights[39][202] = 16'sd-40;
        fc1_weights[39][203] = 16'sd-57;
        fc1_weights[39][204] = 16'sd-57;
        fc1_weights[39][205] = 16'sd-50;
        fc1_weights[39][206] = 16'sd-24;
        fc1_weights[39][207] = 16'sd-1;
        fc1_weights[40][0] = 16'sd2;
        fc1_weights[40][1] = 16'sd5;
        fc1_weights[40][2] = 16'sd-7;
        fc1_weights[40][3] = 16'sd40;
        fc1_weights[40][4] = 16'sd45;
        fc1_weights[40][5] = 16'sd50;
        fc1_weights[40][6] = 16'sd52;
        fc1_weights[40][7] = 16'sd21;
        fc1_weights[40][8] = 16'sd61;
        fc1_weights[40][9] = 16'sd74;
        fc1_weights[40][10] = 16'sd45;
        fc1_weights[40][11] = 16'sd-45;
        fc1_weights[40][12] = 16'sd-21;
        fc1_weights[40][13] = 16'sd-7;
        fc1_weights[40][14] = 16'sd53;
        fc1_weights[40][15] = 16'sd62;
        fc1_weights[40][16] = 16'sd14;
        fc1_weights[40][17] = 16'sd4;
        fc1_weights[40][18] = 16'sd-6;
        fc1_weights[40][19] = 16'sd9;
        fc1_weights[40][20] = 16'sd-3;
        fc1_weights[40][21] = 16'sd11;
        fc1_weights[40][22] = 16'sd70;
        fc1_weights[40][23] = 16'sd14;
        fc1_weights[40][24] = 16'sd30;
        fc1_weights[40][25] = 16'sd13;
        fc1_weights[40][26] = 16'sd-27;
        fc1_weights[40][27] = 16'sd11;
        fc1_weights[40][28] = 16'sd-13;
        fc1_weights[40][29] = 16'sd-6;
        fc1_weights[40][30] = 16'sd22;
        fc1_weights[40][31] = 16'sd19;
        fc1_weights[40][32] = 16'sd18;
        fc1_weights[40][33] = 16'sd18;
        fc1_weights[40][34] = 16'sd20;
        fc1_weights[40][35] = 16'sd60;
        fc1_weights[40][36] = 16'sd67;
        fc1_weights[40][37] = 16'sd35;
        fc1_weights[40][38] = 16'sd-21;
        fc1_weights[40][39] = 16'sd81;
        fc1_weights[40][40] = 16'sd19;
        fc1_weights[40][41] = 16'sd23;
        fc1_weights[40][42] = 16'sd-3;
        fc1_weights[40][43] = 16'sd23;
        fc1_weights[40][44] = 16'sd-17;
        fc1_weights[40][45] = 16'sd-13;
        fc1_weights[40][46] = 16'sd-36;
        fc1_weights[40][47] = 16'sd-9;
        fc1_weights[40][48] = 16'sd32;
        fc1_weights[40][49] = 16'sd32;
        fc1_weights[40][50] = 16'sd-2;
        fc1_weights[40][51] = 16'sd17;
        fc1_weights[40][52] = 16'sd-24;
        fc1_weights[40][53] = 16'sd-16;
        fc1_weights[40][54] = 16'sd-17;
        fc1_weights[40][55] = 16'sd-21;
        fc1_weights[40][56] = 16'sd32;
        fc1_weights[40][57] = 16'sd-2;
        fc1_weights[40][58] = 16'sd-34;
        fc1_weights[40][59] = 16'sd-18;
        fc1_weights[40][60] = 16'sd-9;
        fc1_weights[40][61] = 16'sd-2;
        fc1_weights[40][62] = 16'sd1;
        fc1_weights[40][63] = 16'sd11;
        fc1_weights[40][64] = 16'sd5;
        fc1_weights[40][65] = 16'sd53;
        fc1_weights[40][66] = 16'sd31;
        fc1_weights[40][67] = 16'sd9;
        fc1_weights[40][68] = 16'sd50;
        fc1_weights[40][69] = 16'sd-53;
        fc1_weights[40][70] = 16'sd-25;
        fc1_weights[40][71] = 16'sd32;
        fc1_weights[40][72] = 16'sd-3;
        fc1_weights[40][73] = 16'sd14;
        fc1_weights[40][74] = 16'sd-18;
        fc1_weights[40][75] = 16'sd11;
        fc1_weights[40][76] = 16'sd-12;
        fc1_weights[40][77] = 16'sd-50;
        fc1_weights[40][78] = 16'sd10;
        fc1_weights[40][79] = 16'sd32;
        fc1_weights[40][80] = 16'sd62;
        fc1_weights[40][81] = 16'sd-13;
        fc1_weights[40][82] = 16'sd6;
        fc1_weights[40][83] = 16'sd31;
        fc1_weights[40][84] = 16'sd-22;
        fc1_weights[40][85] = 16'sd-4;
        fc1_weights[40][86] = 16'sd-57;
        fc1_weights[40][87] = 16'sd-11;
        fc1_weights[40][88] = 16'sd-52;
        fc1_weights[40][89] = 16'sd34;
        fc1_weights[40][90] = 16'sd47;
        fc1_weights[40][91] = 16'sd-22;
        fc1_weights[40][92] = 16'sd-52;
        fc1_weights[40][93] = 16'sd29;
        fc1_weights[40][94] = 16'sd0;
        fc1_weights[40][95] = 16'sd11;
        fc1_weights[40][96] = 16'sd-27;
        fc1_weights[40][97] = 16'sd-12;
        fc1_weights[40][98] = 16'sd-27;
        fc1_weights[40][99] = 16'sd55;
        fc1_weights[40][100] = 16'sd-5;
        fc1_weights[40][101] = 16'sd-22;
        fc1_weights[40][102] = 16'sd-35;
        fc1_weights[40][103] = 16'sd-35;
        fc1_weights[40][104] = 16'sd-41;
        fc1_weights[40][105] = 16'sd0;
        fc1_weights[40][106] = 16'sd-39;
        fc1_weights[40][107] = 16'sd-1;
        fc1_weights[40][108] = 16'sd32;
        fc1_weights[40][109] = 16'sd17;
        fc1_weights[40][110] = 16'sd15;
        fc1_weights[40][111] = 16'sd18;
        fc1_weights[40][112] = 16'sd-36;
        fc1_weights[40][113] = 16'sd-33;
        fc1_weights[40][114] = 16'sd-53;
        fc1_weights[40][115] = 16'sd-70;
        fc1_weights[40][116] = 16'sd-21;
        fc1_weights[40][117] = 16'sd16;
        fc1_weights[40][118] = 16'sd5;
        fc1_weights[40][119] = 16'sd14;
        fc1_weights[40][120] = 16'sd17;
        fc1_weights[40][121] = 16'sd20;
        fc1_weights[40][122] = 16'sd11;
        fc1_weights[40][123] = 16'sd7;
        fc1_weights[40][124] = 16'sd42;
        fc1_weights[40][125] = 16'sd40;
        fc1_weights[40][126] = 16'sd21;
        fc1_weights[40][127] = 16'sd17;
        fc1_weights[40][128] = 16'sd-34;
        fc1_weights[40][129] = 16'sd-9;
        fc1_weights[40][130] = 16'sd14;
        fc1_weights[40][131] = 16'sd31;
        fc1_weights[40][132] = 16'sd8;
        fc1_weights[40][133] = 16'sd6;
        fc1_weights[40][134] = 16'sd1;
        fc1_weights[40][135] = 16'sd-28;
        fc1_weights[40][136] = 16'sd-45;
        fc1_weights[40][137] = 16'sd-73;
        fc1_weights[40][138] = 16'sd-107;
        fc1_weights[40][139] = 16'sd-55;
        fc1_weights[40][140] = 16'sd-36;
        fc1_weights[40][141] = 16'sd-61;
        fc1_weights[40][142] = 16'sd15;
        fc1_weights[40][143] = 16'sd52;
        fc1_weights[40][144] = 16'sd-67;
        fc1_weights[40][145] = 16'sd-12;
        fc1_weights[40][146] = 16'sd5;
        fc1_weights[40][147] = 16'sd-14;
        fc1_weights[40][148] = 16'sd-15;
        fc1_weights[40][149] = 16'sd-23;
        fc1_weights[40][150] = 16'sd-30;
        fc1_weights[40][151] = 16'sd-8;
        fc1_weights[40][152] = 16'sd-15;
        fc1_weights[40][153] = 16'sd-31;
        fc1_weights[40][154] = 16'sd-98;
        fc1_weights[40][155] = 16'sd-15;
        fc1_weights[40][156] = 16'sd-11;
        fc1_weights[40][157] = 16'sd-7;
        fc1_weights[40][158] = 16'sd-22;
        fc1_weights[40][159] = 16'sd-54;
        fc1_weights[40][160] = 16'sd-55;
        fc1_weights[40][161] = 16'sd-58;
        fc1_weights[40][162] = 16'sd-51;
        fc1_weights[40][163] = 16'sd-47;
        fc1_weights[40][164] = 16'sd-22;
        fc1_weights[40][165] = 16'sd13;
        fc1_weights[40][166] = 16'sd86;
        fc1_weights[40][167] = 16'sd63;
        fc1_weights[40][168] = 16'sd50;
        fc1_weights[40][169] = 16'sd61;
        fc1_weights[40][170] = 16'sd-4;
        fc1_weights[40][171] = 16'sd-12;
        fc1_weights[40][172] = 16'sd7;
        fc1_weights[40][173] = 16'sd44;
        fc1_weights[40][174] = 16'sd-1;
        fc1_weights[40][175] = 16'sd13;
        fc1_weights[40][176] = 16'sd12;
        fc1_weights[40][177] = 16'sd-18;
        fc1_weights[40][178] = 16'sd-16;
        fc1_weights[40][179] = 16'sd-8;
        fc1_weights[40][180] = 16'sd-79;
        fc1_weights[40][181] = 16'sd-67;
        fc1_weights[40][182] = 16'sd-61;
        fc1_weights[40][183] = 16'sd-36;
        fc1_weights[40][184] = 16'sd-21;
        fc1_weights[40][185] = 16'sd-66;
        fc1_weights[40][186] = 16'sd-38;
        fc1_weights[40][187] = 16'sd-43;
        fc1_weights[40][188] = 16'sd-36;
        fc1_weights[40][189] = 16'sd-27;
        fc1_weights[40][190] = 16'sd-88;
        fc1_weights[40][191] = 16'sd39;
        fc1_weights[40][192] = 16'sd-1;
        fc1_weights[40][193] = 16'sd6;
        fc1_weights[40][194] = 16'sd4;
        fc1_weights[40][195] = 16'sd14;
        fc1_weights[40][196] = 16'sd27;
        fc1_weights[40][197] = 16'sd36;
        fc1_weights[40][198] = 16'sd-11;
        fc1_weights[40][199] = 16'sd8;
        fc1_weights[40][200] = 16'sd-11;
        fc1_weights[40][201] = 16'sd1;
        fc1_weights[40][202] = 16'sd38;
        fc1_weights[40][203] = 16'sd-30;
        fc1_weights[40][204] = 16'sd0;
        fc1_weights[40][205] = 16'sd-11;
        fc1_weights[40][206] = 16'sd-44;
        fc1_weights[40][207] = 16'sd-63;
        fc1_weights[41][0] = 16'sd-10;
        fc1_weights[41][1] = 16'sd20;
        fc1_weights[41][2] = 16'sd50;
        fc1_weights[41][3] = 16'sd-51;
        fc1_weights[41][4] = 16'sd-33;
        fc1_weights[41][5] = 16'sd-9;
        fc1_weights[41][6] = 16'sd-22;
        fc1_weights[41][7] = 16'sd50;
        fc1_weights[41][8] = 16'sd-56;
        fc1_weights[41][9] = 16'sd-100;
        fc1_weights[41][10] = 16'sd27;
        fc1_weights[41][11] = 16'sd-13;
        fc1_weights[41][12] = 16'sd-15;
        fc1_weights[41][13] = 16'sd-20;
        fc1_weights[41][14] = 16'sd-30;
        fc1_weights[41][15] = 16'sd13;
        fc1_weights[41][16] = 16'sd-6;
        fc1_weights[41][17] = 16'sd23;
        fc1_weights[41][18] = 16'sd66;
        fc1_weights[41][19] = 16'sd20;
        fc1_weights[41][20] = 16'sd22;
        fc1_weights[41][21] = 16'sd26;
        fc1_weights[41][22] = 16'sd-7;
        fc1_weights[41][23] = 16'sd20;
        fc1_weights[41][24] = 16'sd45;
        fc1_weights[41][25] = 16'sd65;
        fc1_weights[41][26] = 16'sd3;
        fc1_weights[41][27] = 16'sd-45;
        fc1_weights[41][28] = 16'sd-52;
        fc1_weights[41][29] = 16'sd-6;
        fc1_weights[41][30] = 16'sd29;
        fc1_weights[41][31] = 16'sd-14;
        fc1_weights[41][32] = 16'sd-1;
        fc1_weights[41][33] = 16'sd-13;
        fc1_weights[41][34] = 16'sd-30;
        fc1_weights[41][35] = 16'sd-53;
        fc1_weights[41][36] = 16'sd42;
        fc1_weights[41][37] = 16'sd31;
        fc1_weights[41][38] = 16'sd14;
        fc1_weights[41][39] = 16'sd6;
        fc1_weights[41][40] = 16'sd6;
        fc1_weights[41][41] = 16'sd25;
        fc1_weights[41][42] = 16'sd-10;
        fc1_weights[41][43] = 16'sd39;
        fc1_weights[41][44] = 16'sd24;
        fc1_weights[41][45] = 16'sd-5;
        fc1_weights[41][46] = 16'sd-1;
        fc1_weights[41][47] = 16'sd1;
        fc1_weights[41][48] = 16'sd17;
        fc1_weights[41][49] = 16'sd26;
        fc1_weights[41][50] = 16'sd43;
        fc1_weights[41][51] = 16'sd-12;
        fc1_weights[41][52] = 16'sd-11;
        fc1_weights[41][53] = 16'sd24;
        fc1_weights[41][54] = 16'sd-40;
        fc1_weights[41][55] = 16'sd75;
        fc1_weights[41][56] = 16'sd10;
        fc1_weights[41][57] = 16'sd33;
        fc1_weights[41][58] = 16'sd25;
        fc1_weights[41][59] = 16'sd4;
        fc1_weights[41][60] = 16'sd-10;
        fc1_weights[41][61] = 16'sd25;
        fc1_weights[41][62] = 16'sd-11;
        fc1_weights[41][63] = 16'sd23;
        fc1_weights[41][64] = 16'sd69;
        fc1_weights[41][65] = 16'sd-43;
        fc1_weights[41][66] = 16'sd-19;
        fc1_weights[41][67] = 16'sd-60;
        fc1_weights[41][68] = 16'sd-23;
        fc1_weights[41][69] = 16'sd39;
        fc1_weights[41][70] = 16'sd46;
        fc1_weights[41][71] = 16'sd-9;
        fc1_weights[41][72] = 16'sd-19;
        fc1_weights[41][73] = 16'sd-1;
        fc1_weights[41][74] = 16'sd-8;
        fc1_weights[41][75] = 16'sd-47;
        fc1_weights[41][76] = 16'sd-47;
        fc1_weights[41][77] = 16'sd11;
        fc1_weights[41][78] = 16'sd-39;
        fc1_weights[41][79] = 16'sd-48;
        fc1_weights[41][80] = 16'sd-25;
        fc1_weights[41][81] = 16'sd-20;
        fc1_weights[41][82] = 16'sd-76;
        fc1_weights[41][83] = 16'sd64;
        fc1_weights[41][84] = 16'sd12;
        fc1_weights[41][85] = 16'sd4;
        fc1_weights[41][86] = 16'sd-38;
        fc1_weights[41][87] = 16'sd-6;
        fc1_weights[41][88] = 16'sd-47;
        fc1_weights[41][89] = 16'sd-28;
        fc1_weights[41][90] = 16'sd-7;
        fc1_weights[41][91] = 16'sd-67;
        fc1_weights[41][92] = 16'sd-51;
        fc1_weights[41][93] = 16'sd-32;
        fc1_weights[41][94] = 16'sd-89;
        fc1_weights[41][95] = 16'sd-41;
        fc1_weights[41][96] = 16'sd-20;
        fc1_weights[41][97] = 16'sd18;
        fc1_weights[41][98] = 16'sd-7;
        fc1_weights[41][99] = 16'sd-2;
        fc1_weights[41][100] = 16'sd-30;
        fc1_weights[41][101] = 16'sd-47;
        fc1_weights[41][102] = 16'sd-76;
        fc1_weights[41][103] = 16'sd-56;
        fc1_weights[41][104] = 16'sd-28;
        fc1_weights[41][105] = 16'sd-28;
        fc1_weights[41][106] = 16'sd12;
        fc1_weights[41][107] = 16'sd-59;
        fc1_weights[41][108] = 16'sd18;
        fc1_weights[41][109] = 16'sd33;
        fc1_weights[41][110] = 16'sd40;
        fc1_weights[41][111] = 16'sd15;
        fc1_weights[41][112] = 16'sd25;
        fc1_weights[41][113] = 16'sd44;
        fc1_weights[41][114] = 16'sd41;
        fc1_weights[41][115] = 16'sd93;
        fc1_weights[41][116] = 16'sd-18;
        fc1_weights[41][117] = 16'sd13;
        fc1_weights[41][118] = 16'sd-24;
        fc1_weights[41][119] = 16'sd-74;
        fc1_weights[41][120] = 16'sd-94;
        fc1_weights[41][121] = 16'sd-40;
        fc1_weights[41][122] = 16'sd-24;
        fc1_weights[41][123] = 16'sd-25;
        fc1_weights[41][124] = 16'sd-96;
        fc1_weights[41][125] = 16'sd-67;
        fc1_weights[41][126] = 16'sd-15;
        fc1_weights[41][127] = 16'sd35;
        fc1_weights[41][128] = 16'sd-51;
        fc1_weights[41][129] = 16'sd-50;
        fc1_weights[41][130] = 16'sd15;
        fc1_weights[41][131] = 16'sd4;
        fc1_weights[41][132] = 16'sd14;
        fc1_weights[41][133] = 16'sd-3;
        fc1_weights[41][134] = 16'sd16;
        fc1_weights[41][135] = 16'sd4;
        fc1_weights[41][136] = 16'sd63;
        fc1_weights[41][137] = 16'sd-19;
        fc1_weights[41][138] = 16'sd116;
        fc1_weights[41][139] = 16'sd-37;
        fc1_weights[41][140] = 16'sd-46;
        fc1_weights[41][141] = 16'sd25;
        fc1_weights[41][142] = 16'sd-62;
        fc1_weights[41][143] = 16'sd39;
        fc1_weights[41][144] = 16'sd18;
        fc1_weights[41][145] = 16'sd10;
        fc1_weights[41][146] = 16'sd29;
        fc1_weights[41][147] = 16'sd49;
        fc1_weights[41][148] = 16'sd14;
        fc1_weights[41][149] = 16'sd-11;
        fc1_weights[41][150] = 16'sd6;
        fc1_weights[41][151] = 16'sd27;
        fc1_weights[41][152] = 16'sd20;
        fc1_weights[41][153] = 16'sd-32;
        fc1_weights[41][154] = 16'sd-29;
        fc1_weights[41][155] = 16'sd-5;
        fc1_weights[41][156] = 16'sd-36;
        fc1_weights[41][157] = 16'sd-31;
        fc1_weights[41][158] = 16'sd13;
        fc1_weights[41][159] = 16'sd29;
        fc1_weights[41][160] = 16'sd54;
        fc1_weights[41][161] = 16'sd35;
        fc1_weights[41][162] = 16'sd44;
        fc1_weights[41][163] = 16'sd-32;
        fc1_weights[41][164] = 16'sd1;
        fc1_weights[41][165] = 16'sd-11;
        fc1_weights[41][166] = 16'sd5;
        fc1_weights[41][167] = 16'sd17;
        fc1_weights[41][168] = 16'sd-13;
        fc1_weights[41][169] = 16'sd8;
        fc1_weights[41][170] = 16'sd63;
        fc1_weights[41][171] = 16'sd-27;
        fc1_weights[41][172] = 16'sd72;
        fc1_weights[41][173] = 16'sd1;
        fc1_weights[41][174] = 16'sd-12;
        fc1_weights[41][175] = 16'sd10;
        fc1_weights[41][176] = 16'sd59;
        fc1_weights[41][177] = 16'sd76;
        fc1_weights[41][178] = 16'sd-23;
        fc1_weights[41][179] = 16'sd13;
        fc1_weights[41][180] = 16'sd2;
        fc1_weights[41][181] = 16'sd17;
        fc1_weights[41][182] = 16'sd-22;
        fc1_weights[41][183] = 16'sd-33;
        fc1_weights[41][184] = 16'sd-33;
        fc1_weights[41][185] = 16'sd2;
        fc1_weights[41][186] = 16'sd31;
        fc1_weights[41][187] = 16'sd-11;
        fc1_weights[41][188] = 16'sd-18;
        fc1_weights[41][189] = 16'sd-28;
        fc1_weights[41][190] = 16'sd-12;
        fc1_weights[41][191] = 16'sd-6;
        fc1_weights[41][192] = 16'sd-25;
        fc1_weights[41][193] = 16'sd-21;
        fc1_weights[41][194] = 16'sd-72;
        fc1_weights[41][195] = 16'sd15;
        fc1_weights[41][196] = 16'sd55;
        fc1_weights[41][197] = 16'sd40;
        fc1_weights[41][198] = 16'sd9;
        fc1_weights[41][199] = 16'sd57;
        fc1_weights[41][200] = 16'sd58;
        fc1_weights[41][201] = 16'sd7;
        fc1_weights[41][202] = 16'sd-1;
        fc1_weights[41][203] = 16'sd69;
        fc1_weights[41][204] = 16'sd110;
        fc1_weights[41][205] = 16'sd84;
        fc1_weights[41][206] = 16'sd25;
        fc1_weights[41][207] = 16'sd11;
        fc1_weights[42][0] = 16'sd-107;
        fc1_weights[42][1] = 16'sd-49;
        fc1_weights[42][2] = 16'sd-14;
        fc1_weights[42][3] = 16'sd-64;
        fc1_weights[42][4] = 16'sd-38;
        fc1_weights[42][5] = 16'sd-22;
        fc1_weights[42][6] = 16'sd-13;
        fc1_weights[42][7] = 16'sd-6;
        fc1_weights[42][8] = 16'sd17;
        fc1_weights[42][9] = 16'sd-1;
        fc1_weights[42][10] = 16'sd17;
        fc1_weights[42][11] = 16'sd33;
        fc1_weights[42][12] = 16'sd29;
        fc1_weights[42][13] = 16'sd28;
        fc1_weights[42][14] = 16'sd13;
        fc1_weights[42][15] = 16'sd13;
        fc1_weights[42][16] = 16'sd10;
        fc1_weights[42][17] = 16'sd21;
        fc1_weights[42][18] = 16'sd5;
        fc1_weights[42][19] = 16'sd-9;
        fc1_weights[42][20] = 16'sd-35;
        fc1_weights[42][21] = 16'sd18;
        fc1_weights[42][22] = 16'sd21;
        fc1_weights[42][23] = 16'sd18;
        fc1_weights[42][24] = 16'sd-21;
        fc1_weights[42][25] = 16'sd-11;
        fc1_weights[42][26] = 16'sd-43;
        fc1_weights[42][27] = 16'sd-54;
        fc1_weights[42][28] = 16'sd-27;
        fc1_weights[42][29] = 16'sd-42;
        fc1_weights[42][30] = 16'sd-15;
        fc1_weights[42][31] = 16'sd4;
        fc1_weights[42][32] = 16'sd3;
        fc1_weights[42][33] = 16'sd-24;
        fc1_weights[42][34] = 16'sd-36;
        fc1_weights[42][35] = 16'sd-54;
        fc1_weights[42][36] = 16'sd0;
        fc1_weights[42][37] = 16'sd43;
        fc1_weights[42][38] = 16'sd-26;
        fc1_weights[42][39] = 16'sd29;
        fc1_weights[42][40] = 16'sd-28;
        fc1_weights[42][41] = 16'sd-21;
        fc1_weights[42][42] = 16'sd20;
        fc1_weights[42][43] = 16'sd8;
        fc1_weights[42][44] = 16'sd-6;
        fc1_weights[42][45] = 16'sd-24;
        fc1_weights[42][46] = 16'sd-42;
        fc1_weights[42][47] = 16'sd-22;
        fc1_weights[42][48] = 16'sd-20;
        fc1_weights[42][49] = 16'sd-9;
        fc1_weights[42][50] = 16'sd13;
        fc1_weights[42][51] = 16'sd-16;
        fc1_weights[42][52] = 16'sd4;
        fc1_weights[42][53] = 16'sd-20;
        fc1_weights[42][54] = 16'sd-42;
        fc1_weights[42][55] = 16'sd-30;
        fc1_weights[42][56] = 16'sd22;
        fc1_weights[42][57] = 16'sd0;
        fc1_weights[42][58] = 16'sd-16;
        fc1_weights[42][59] = 16'sd-7;
        fc1_weights[42][60] = 16'sd-18;
        fc1_weights[42][61] = 16'sd-40;
        fc1_weights[42][62] = 16'sd-30;
        fc1_weights[42][63] = 16'sd-1;
        fc1_weights[42][64] = 16'sd-26;
        fc1_weights[42][65] = 16'sd-6;
        fc1_weights[42][66] = 16'sd27;
        fc1_weights[42][67] = 16'sd-29;
        fc1_weights[42][68] = 16'sd8;
        fc1_weights[42][69] = 16'sd16;
        fc1_weights[42][70] = 16'sd6;
        fc1_weights[42][71] = 16'sd-42;
        fc1_weights[42][72] = 16'sd-43;
        fc1_weights[42][73] = 16'sd15;
        fc1_weights[42][74] = 16'sd-20;
        fc1_weights[42][75] = 16'sd18;
        fc1_weights[42][76] = 16'sd8;
        fc1_weights[42][77] = 16'sd-3;
        fc1_weights[42][78] = 16'sd-37;
        fc1_weights[42][79] = 16'sd-34;
        fc1_weights[42][80] = 16'sd-10;
        fc1_weights[42][81] = 16'sd-10;
        fc1_weights[42][82] = 16'sd-13;
        fc1_weights[42][83] = 16'sd12;
        fc1_weights[42][84] = 16'sd-3;
        fc1_weights[42][85] = 16'sd22;
        fc1_weights[42][86] = 16'sd35;
        fc1_weights[42][87] = 16'sd16;
        fc1_weights[42][88] = 16'sd5;
        fc1_weights[42][89] = 16'sd-17;
        fc1_weights[42][90] = 16'sd1;
        fc1_weights[42][91] = 16'sd-6;
        fc1_weights[42][92] = 16'sd10;
        fc1_weights[42][93] = 16'sd-40;
        fc1_weights[42][94] = 16'sd-16;
        fc1_weights[42][95] = 16'sd10;
        fc1_weights[42][96] = 16'sd-18;
        fc1_weights[42][97] = 16'sd-26;
        fc1_weights[42][98] = 16'sd7;
        fc1_weights[42][99] = 16'sd12;
        fc1_weights[42][100] = 16'sd-18;
        fc1_weights[42][101] = 16'sd12;
        fc1_weights[42][102] = 16'sd-2;
        fc1_weights[42][103] = 16'sd10;
        fc1_weights[42][104] = 16'sd-10;
        fc1_weights[42][105] = 16'sd18;
        fc1_weights[42][106] = 16'sd28;
        fc1_weights[42][107] = 16'sd-1;
        fc1_weights[42][108] = 16'sd5;
        fc1_weights[42][109] = 16'sd29;
        fc1_weights[42][110] = 16'sd53;
        fc1_weights[42][111] = 16'sd73;
        fc1_weights[42][112] = 16'sd33;
        fc1_weights[42][113] = 16'sd-15;
        fc1_weights[42][114] = 16'sd34;
        fc1_weights[42][115] = 16'sd56;
        fc1_weights[42][116] = 16'sd-40;
        fc1_weights[42][117] = 16'sd-28;
        fc1_weights[42][118] = 16'sd0;
        fc1_weights[42][119] = 16'sd-5;
        fc1_weights[42][120] = 16'sd-12;
        fc1_weights[42][121] = 16'sd-2;
        fc1_weights[42][122] = 16'sd-19;
        fc1_weights[42][123] = 16'sd-11;
        fc1_weights[42][124] = 16'sd-9;
        fc1_weights[42][125] = 16'sd-5;
        fc1_weights[42][126] = 16'sd-13;
        fc1_weights[42][127] = 16'sd31;
        fc1_weights[42][128] = 16'sd31;
        fc1_weights[42][129] = 16'sd38;
        fc1_weights[42][130] = 16'sd4;
        fc1_weights[42][131] = 16'sd10;
        fc1_weights[42][132] = 16'sd9;
        fc1_weights[42][133] = 16'sd7;
        fc1_weights[42][134] = 16'sd-9;
        fc1_weights[42][135] = 16'sd3;
        fc1_weights[42][136] = 16'sd-3;
        fc1_weights[42][137] = 16'sd2;
        fc1_weights[42][138] = 16'sd3;
        fc1_weights[42][139] = 16'sd24;
        fc1_weights[42][140] = 16'sd55;
        fc1_weights[42][141] = 16'sd85;
        fc1_weights[42][142] = 16'sd2;
        fc1_weights[42][143] = 16'sd26;
        fc1_weights[42][144] = 16'sd-12;
        fc1_weights[42][145] = 16'sd2;
        fc1_weights[42][146] = 16'sd-25;
        fc1_weights[42][147] = 16'sd-56;
        fc1_weights[42][148] = 16'sd-20;
        fc1_weights[42][149] = 16'sd-32;
        fc1_weights[42][150] = 16'sd8;
        fc1_weights[42][151] = 16'sd-24;
        fc1_weights[42][152] = 16'sd0;
        fc1_weights[42][153] = 16'sd-2;
        fc1_weights[42][154] = 16'sd0;
        fc1_weights[42][155] = 16'sd-27;
        fc1_weights[42][156] = 16'sd15;
        fc1_weights[42][157] = 16'sd25;
        fc1_weights[42][158] = 16'sd7;
        fc1_weights[42][159] = 16'sd-25;
        fc1_weights[42][160] = 16'sd29;
        fc1_weights[42][161] = 16'sd23;
        fc1_weights[42][162] = 16'sd27;
        fc1_weights[42][163] = 16'sd12;
        fc1_weights[42][164] = 16'sd34;
        fc1_weights[42][165] = 16'sd5;
        fc1_weights[42][166] = 16'sd4;
        fc1_weights[42][167] = 16'sd12;
        fc1_weights[42][168] = 16'sd11;
        fc1_weights[42][169] = 16'sd-2;
        fc1_weights[42][170] = 16'sd5;
        fc1_weights[42][171] = 16'sd-25;
        fc1_weights[42][172] = 16'sd-18;
        fc1_weights[42][173] = 16'sd-8;
        fc1_weights[42][174] = 16'sd-10;
        fc1_weights[42][175] = 16'sd-39;
        fc1_weights[42][176] = 16'sd-15;
        fc1_weights[42][177] = 16'sd-10;
        fc1_weights[42][178] = 16'sd-30;
        fc1_weights[42][179] = 16'sd-9;
        fc1_weights[42][180] = 16'sd-46;
        fc1_weights[42][181] = 16'sd-49;
        fc1_weights[42][182] = 16'sd38;
        fc1_weights[42][183] = 16'sd22;
        fc1_weights[42][184] = 16'sd13;
        fc1_weights[42][185] = 16'sd-15;
        fc1_weights[42][186] = 16'sd25;
        fc1_weights[42][187] = 16'sd9;
        fc1_weights[42][188] = 16'sd7;
        fc1_weights[42][189] = 16'sd8;
        fc1_weights[42][190] = 16'sd5;
        fc1_weights[42][191] = 16'sd28;
        fc1_weights[42][192] = 16'sd32;
        fc1_weights[42][193] = 16'sd30;
        fc1_weights[42][194] = 16'sd3;
        fc1_weights[42][195] = 16'sd16;
        fc1_weights[42][196] = 16'sd6;
        fc1_weights[42][197] = 16'sd-12;
        fc1_weights[42][198] = 16'sd-15;
        fc1_weights[42][199] = 16'sd5;
        fc1_weights[42][200] = 16'sd-16;
        fc1_weights[42][201] = 16'sd-19;
        fc1_weights[42][202] = 16'sd-18;
        fc1_weights[42][203] = 16'sd-29;
        fc1_weights[42][204] = 16'sd-10;
        fc1_weights[42][205] = 16'sd-24;
        fc1_weights[42][206] = 16'sd9;
        fc1_weights[42][207] = 16'sd6;
        fc1_weights[43][0] = 16'sd15;
        fc1_weights[43][1] = 16'sd-2;
        fc1_weights[43][2] = 16'sd40;
        fc1_weights[43][3] = 16'sd24;
        fc1_weights[43][4] = 16'sd-49;
        fc1_weights[43][5] = 16'sd-11;
        fc1_weights[43][6] = 16'sd17;
        fc1_weights[43][7] = 16'sd-16;
        fc1_weights[43][8] = 16'sd-30;
        fc1_weights[43][9] = 16'sd-5;
        fc1_weights[43][10] = 16'sd17;
        fc1_weights[43][11] = 16'sd23;
        fc1_weights[43][12] = 16'sd83;
        fc1_weights[43][13] = 16'sd61;
        fc1_weights[43][14] = 16'sd57;
        fc1_weights[43][15] = 16'sd-19;
        fc1_weights[43][16] = 16'sd-22;
        fc1_weights[43][17] = 16'sd23;
        fc1_weights[43][18] = 16'sd16;
        fc1_weights[43][19] = 16'sd36;
        fc1_weights[43][20] = 16'sd-31;
        fc1_weights[43][21] = 16'sd-12;
        fc1_weights[43][22] = 16'sd-20;
        fc1_weights[43][23] = 16'sd-11;
        fc1_weights[43][24] = 16'sd-6;
        fc1_weights[43][25] = 16'sd-12;
        fc1_weights[43][26] = 16'sd48;
        fc1_weights[43][27] = 16'sd-1;
        fc1_weights[43][28] = 16'sd14;
        fc1_weights[43][29] = 16'sd7;
        fc1_weights[43][30] = 16'sd-17;
        fc1_weights[43][31] = 16'sd-24;
        fc1_weights[43][32] = 16'sd-12;
        fc1_weights[43][33] = 16'sd32;
        fc1_weights[43][34] = 16'sd-19;
        fc1_weights[43][35] = 16'sd4;
        fc1_weights[43][36] = 16'sd-15;
        fc1_weights[43][37] = 16'sd43;
        fc1_weights[43][38] = 16'sd81;
        fc1_weights[43][39] = 16'sd31;
        fc1_weights[43][40] = 16'sd29;
        fc1_weights[43][41] = 16'sd-8;
        fc1_weights[43][42] = 16'sd-16;
        fc1_weights[43][43] = 16'sd1;
        fc1_weights[43][44] = 16'sd35;
        fc1_weights[43][45] = 16'sd23;
        fc1_weights[43][46] = 16'sd37;
        fc1_weights[43][47] = 16'sd25;
        fc1_weights[43][48] = 16'sd27;
        fc1_weights[43][49] = 16'sd-42;
        fc1_weights[43][50] = 16'sd4;
        fc1_weights[43][51] = 16'sd-24;
        fc1_weights[43][52] = 16'sd20;
        fc1_weights[43][53] = 16'sd34;
        fc1_weights[43][54] = 16'sd11;
        fc1_weights[43][55] = 16'sd-4;
        fc1_weights[43][56] = 16'sd-43;
        fc1_weights[43][57] = 16'sd-3;
        fc1_weights[43][58] = 16'sd-1;
        fc1_weights[43][59] = 16'sd2;
        fc1_weights[43][60] = 16'sd-6;
        fc1_weights[43][61] = 16'sd10;
        fc1_weights[43][62] = 16'sd-1;
        fc1_weights[43][63] = 16'sd22;
        fc1_weights[43][64] = 16'sd20;
        fc1_weights[43][65] = 16'sd66;
        fc1_weights[43][66] = 16'sd-19;
        fc1_weights[43][67] = 16'sd-7;
        fc1_weights[43][68] = 16'sd8;
        fc1_weights[43][69] = 16'sd6;
        fc1_weights[43][70] = 16'sd3;
        fc1_weights[43][71] = 16'sd-24;
        fc1_weights[43][72] = 16'sd-13;
        fc1_weights[43][73] = 16'sd18;
        fc1_weights[43][74] = 16'sd-14;
        fc1_weights[43][75] = 16'sd-12;
        fc1_weights[43][76] = 16'sd-35;
        fc1_weights[43][77] = 16'sd-29;
        fc1_weights[43][78] = 16'sd30;
        fc1_weights[43][79] = 16'sd-51;
        fc1_weights[43][80] = 16'sd-46;
        fc1_weights[43][81] = 16'sd-30;
        fc1_weights[43][82] = 16'sd-20;
        fc1_weights[43][83] = 16'sd-56;
        fc1_weights[43][84] = 16'sd0;
        fc1_weights[43][85] = 16'sd54;
        fc1_weights[43][86] = 16'sd14;
        fc1_weights[43][87] = 16'sd-16;
        fc1_weights[43][88] = 16'sd6;
        fc1_weights[43][89] = 16'sd27;
        fc1_weights[43][90] = 16'sd-56;
        fc1_weights[43][91] = 16'sd-16;
        fc1_weights[43][92] = 16'sd-28;
        fc1_weights[43][93] = 16'sd-27;
        fc1_weights[43][94] = 16'sd29;
        fc1_weights[43][95] = 16'sd-17;
        fc1_weights[43][96] = 16'sd50;
        fc1_weights[43][97] = 16'sd-6;
        fc1_weights[43][98] = 16'sd13;
        fc1_weights[43][99] = 16'sd6;
        fc1_weights[43][100] = 16'sd-38;
        fc1_weights[43][101] = 16'sd17;
        fc1_weights[43][102] = 16'sd-4;
        fc1_weights[43][103] = 16'sd13;
        fc1_weights[43][104] = 16'sd-4;
        fc1_weights[43][105] = 16'sd30;
        fc1_weights[43][106] = 16'sd11;
        fc1_weights[43][107] = 16'sd-30;
        fc1_weights[43][108] = 16'sd-21;
        fc1_weights[43][109] = 16'sd-39;
        fc1_weights[43][110] = 16'sd-1;
        fc1_weights[43][111] = 16'sd-34;
        fc1_weights[43][112] = 16'sd-105;
        fc1_weights[43][113] = 16'sd-62;
        fc1_weights[43][114] = 16'sd21;
        fc1_weights[43][115] = 16'sd48;
        fc1_weights[43][116] = 16'sd-12;
        fc1_weights[43][117] = 16'sd-65;
        fc1_weights[43][118] = 16'sd-22;
        fc1_weights[43][119] = 16'sd-44;
        fc1_weights[43][120] = 16'sd-41;
        fc1_weights[43][121] = 16'sd-40;
        fc1_weights[43][122] = 16'sd-16;
        fc1_weights[43][123] = 16'sd-56;
        fc1_weights[43][124] = 16'sd-17;
        fc1_weights[43][125] = 16'sd-31;
        fc1_weights[43][126] = 16'sd-47;
        fc1_weights[43][127] = 16'sd-50;
        fc1_weights[43][128] = 16'sd-43;
        fc1_weights[43][129] = 16'sd-1;
        fc1_weights[43][130] = 16'sd2;
        fc1_weights[43][131] = 16'sd42;
        fc1_weights[43][132] = 16'sd43;
        fc1_weights[43][133] = 16'sd6;
        fc1_weights[43][134] = 16'sd2;
        fc1_weights[43][135] = 16'sd-30;
        fc1_weights[43][136] = 16'sd-31;
        fc1_weights[43][137] = 16'sd-21;
        fc1_weights[43][138] = 16'sd32;
        fc1_weights[43][139] = 16'sd35;
        fc1_weights[43][140] = 16'sd51;
        fc1_weights[43][141] = 16'sd33;
        fc1_weights[43][142] = 16'sd-21;
        fc1_weights[43][143] = 16'sd48;
        fc1_weights[43][144] = 16'sd9;
        fc1_weights[43][145] = 16'sd-9;
        fc1_weights[43][146] = 16'sd-12;
        fc1_weights[43][147] = 16'sd-29;
        fc1_weights[43][148] = 16'sd-18;
        fc1_weights[43][149] = 16'sd-8;
        fc1_weights[43][150] = 16'sd26;
        fc1_weights[43][151] = 16'sd-11;
        fc1_weights[43][152] = 16'sd29;
        fc1_weights[43][153] = 16'sd3;
        fc1_weights[43][154] = 16'sd16;
        fc1_weights[43][155] = 16'sd-18;
        fc1_weights[43][156] = 16'sd-48;
        fc1_weights[43][157] = 16'sd-30;
        fc1_weights[43][158] = 16'sd11;
        fc1_weights[43][159] = 16'sd-28;
        fc1_weights[43][160] = 16'sd52;
        fc1_weights[43][161] = 16'sd4;
        fc1_weights[43][162] = 16'sd-55;
        fc1_weights[43][163] = 16'sd-42;
        fc1_weights[43][164] = 16'sd5;
        fc1_weights[43][165] = 16'sd45;
        fc1_weights[43][166] = 16'sd27;
        fc1_weights[43][167] = 16'sd45;
        fc1_weights[43][168] = 16'sd67;
        fc1_weights[43][169] = 16'sd40;
        fc1_weights[43][170] = 16'sd-1;
        fc1_weights[43][171] = 16'sd-11;
        fc1_weights[43][172] = 16'sd-48;
        fc1_weights[43][173] = 16'sd-7;
        fc1_weights[43][174] = 16'sd-27;
        fc1_weights[43][175] = 16'sd-20;
        fc1_weights[43][176] = 16'sd-18;
        fc1_weights[43][177] = 16'sd-29;
        fc1_weights[43][178] = 16'sd-3;
        fc1_weights[43][179] = 16'sd-10;
        fc1_weights[43][180] = 16'sd15;
        fc1_weights[43][181] = 16'sd42;
        fc1_weights[43][182] = 16'sd32;
        fc1_weights[43][183] = 16'sd32;
        fc1_weights[43][184] = 16'sd34;
        fc1_weights[43][185] = 16'sd1;
        fc1_weights[43][186] = 16'sd-46;
        fc1_weights[43][187] = 16'sd0;
        fc1_weights[43][188] = 16'sd18;
        fc1_weights[43][189] = 16'sd4;
        fc1_weights[43][190] = 16'sd16;
        fc1_weights[43][191] = 16'sd33;
        fc1_weights[43][192] = 16'sd18;
        fc1_weights[43][193] = 16'sd38;
        fc1_weights[43][194] = 16'sd16;
        fc1_weights[43][195] = 16'sd-8;
        fc1_weights[43][196] = 16'sd12;
        fc1_weights[43][197] = 16'sd-39;
        fc1_weights[43][198] = 16'sd20;
        fc1_weights[43][199] = 16'sd-33;
        fc1_weights[43][200] = 16'sd-30;
        fc1_weights[43][201] = 16'sd12;
        fc1_weights[43][202] = 16'sd-32;
        fc1_weights[43][203] = 16'sd-43;
        fc1_weights[43][204] = 16'sd-18;
        fc1_weights[43][205] = 16'sd18;
        fc1_weights[43][206] = 16'sd-3;
        fc1_weights[43][207] = 16'sd1;
        fc1_weights[44][0] = 16'sd72;
        fc1_weights[44][1] = 16'sd47;
        fc1_weights[44][2] = 16'sd-16;
        fc1_weights[44][3] = 16'sd-7;
        fc1_weights[44][4] = 16'sd39;
        fc1_weights[44][5] = 16'sd-37;
        fc1_weights[44][6] = 16'sd-59;
        fc1_weights[44][7] = 16'sd-4;
        fc1_weights[44][8] = 16'sd-7;
        fc1_weights[44][9] = 16'sd12;
        fc1_weights[44][10] = 16'sd-46;
        fc1_weights[44][11] = 16'sd-22;
        fc1_weights[44][12] = 16'sd-1;
        fc1_weights[44][13] = 16'sd-16;
        fc1_weights[44][14] = 16'sd2;
        fc1_weights[44][15] = 16'sd41;
        fc1_weights[44][16] = 16'sd-60;
        fc1_weights[44][17] = 16'sd-18;
        fc1_weights[44][18] = 16'sd-20;
        fc1_weights[44][19] = 16'sd-22;
        fc1_weights[44][20] = 16'sd68;
        fc1_weights[44][21] = 16'sd53;
        fc1_weights[44][22] = 16'sd24;
        fc1_weights[44][23] = 16'sd-28;
        fc1_weights[44][24] = 16'sd68;
        fc1_weights[44][25] = 16'sd35;
        fc1_weights[44][26] = 16'sd31;
        fc1_weights[44][27] = 16'sd33;
        fc1_weights[44][28] = 16'sd45;
        fc1_weights[44][29] = 16'sd9;
        fc1_weights[44][30] = 16'sd31;
        fc1_weights[44][31] = 16'sd-35;
        fc1_weights[44][32] = 16'sd-74;
        fc1_weights[44][33] = 16'sd-48;
        fc1_weights[44][34] = 16'sd-51;
        fc1_weights[44][35] = 16'sd-11;
        fc1_weights[44][36] = 16'sd9;
        fc1_weights[44][37] = 16'sd-85;
        fc1_weights[44][38] = 16'sd12;
        fc1_weights[44][39] = 16'sd20;
        fc1_weights[44][40] = 16'sd34;
        fc1_weights[44][41] = 16'sd22;
        fc1_weights[44][42] = 16'sd-23;
        fc1_weights[44][43] = 16'sd51;
        fc1_weights[44][44] = 16'sd-14;
        fc1_weights[44][45] = 16'sd-1;
        fc1_weights[44][46] = 16'sd6;
        fc1_weights[44][47] = 16'sd106;
        fc1_weights[44][48] = 16'sd12;
        fc1_weights[44][49] = 16'sd-32;
        fc1_weights[44][50] = 16'sd-7;
        fc1_weights[44][51] = 16'sd-35;
        fc1_weights[44][52] = 16'sd-2;
        fc1_weights[44][53] = 16'sd56;
        fc1_weights[44][54] = 16'sd20;
        fc1_weights[44][55] = 16'sd44;
        fc1_weights[44][56] = 16'sd4;
        fc1_weights[44][57] = 16'sd11;
        fc1_weights[44][58] = 16'sd-8;
        fc1_weights[44][59] = 16'sd5;
        fc1_weights[44][60] = 16'sd-41;
        fc1_weights[44][61] = 16'sd8;
        fc1_weights[44][62] = 16'sd-45;
        fc1_weights[44][63] = 16'sd-35;
        fc1_weights[44][64] = 16'sd18;
        fc1_weights[44][65] = 16'sd-67;
        fc1_weights[44][66] = 16'sd-28;
        fc1_weights[44][67] = 16'sd30;
        fc1_weights[44][68] = 16'sd-2;
        fc1_weights[44][69] = 16'sd18;
        fc1_weights[44][70] = 16'sd-4;
        fc1_weights[44][71] = 16'sd56;
        fc1_weights[44][72] = 16'sd79;
        fc1_weights[44][73] = 16'sd39;
        fc1_weights[44][74] = 16'sd-23;
        fc1_weights[44][75] = 16'sd12;
        fc1_weights[44][76] = 16'sd-15;
        fc1_weights[44][77] = 16'sd1;
        fc1_weights[44][78] = 16'sd24;
        fc1_weights[44][79] = 16'sd87;
        fc1_weights[44][80] = 16'sd-21;
        fc1_weights[44][81] = 16'sd-23;
        fc1_weights[44][82] = 16'sd16;
        fc1_weights[44][83] = 16'sd-53;
        fc1_weights[44][84] = 16'sd5;
        fc1_weights[44][85] = 16'sd-13;
        fc1_weights[44][86] = 16'sd21;
        fc1_weights[44][87] = 16'sd-12;
        fc1_weights[44][88] = 16'sd-18;
        fc1_weights[44][89] = 16'sd-38;
        fc1_weights[44][90] = 16'sd45;
        fc1_weights[44][91] = 16'sd39;
        fc1_weights[44][92] = 16'sd22;
        fc1_weights[44][93] = 16'sd-22;
        fc1_weights[44][94] = 16'sd-44;
        fc1_weights[44][95] = 16'sd-5;
        fc1_weights[44][96] = 16'sd-47;
        fc1_weights[44][97] = 16'sd-35;
        fc1_weights[44][98] = 16'sd18;
        fc1_weights[44][99] = 16'sd0;
        fc1_weights[44][100] = 16'sd19;
        fc1_weights[44][101] = 16'sd-11;
        fc1_weights[44][102] = 16'sd0;
        fc1_weights[44][103] = 16'sd-46;
        fc1_weights[44][104] = 16'sd68;
        fc1_weights[44][105] = 16'sd6;
        fc1_weights[44][106] = 16'sd29;
        fc1_weights[44][107] = 16'sd28;
        fc1_weights[44][108] = 16'sd8;
        fc1_weights[44][109] = 16'sd-65;
        fc1_weights[44][110] = 16'sd36;
        fc1_weights[44][111] = 16'sd-24;
        fc1_weights[44][112] = 16'sd21;
        fc1_weights[44][113] = 16'sd55;
        fc1_weights[44][114] = 16'sd6;
        fc1_weights[44][115] = 16'sd-42;
        fc1_weights[44][116] = 16'sd23;
        fc1_weights[44][117] = 16'sd-4;
        fc1_weights[44][118] = 16'sd-21;
        fc1_weights[44][119] = 16'sd-32;
        fc1_weights[44][120] = 16'sd-54;
        fc1_weights[44][121] = 16'sd-21;
        fc1_weights[44][122] = 16'sd-26;
        fc1_weights[44][123] = 16'sd4;
        fc1_weights[44][124] = 16'sd-39;
        fc1_weights[44][125] = 16'sd17;
        fc1_weights[44][126] = 16'sd-66;
        fc1_weights[44][127] = 16'sd-34;
        fc1_weights[44][128] = 16'sd-25;
        fc1_weights[44][129] = 16'sd-128;
        fc1_weights[44][130] = 16'sd45;
        fc1_weights[44][131] = 16'sd-38;
        fc1_weights[44][132] = 16'sd-47;
        fc1_weights[44][133] = 16'sd-43;
        fc1_weights[44][134] = 16'sd-32;
        fc1_weights[44][135] = 16'sd-48;
        fc1_weights[44][136] = 16'sd36;
        fc1_weights[44][137] = 16'sd44;
        fc1_weights[44][138] = 16'sd-19;
        fc1_weights[44][139] = 16'sd-12;
        fc1_weights[44][140] = 16'sd-61;
        fc1_weights[44][141] = 16'sd-75;
        fc1_weights[44][142] = 16'sd-32;
        fc1_weights[44][143] = 16'sd-50;
        fc1_weights[44][144] = 16'sd-66;
        fc1_weights[44][145] = 16'sd-70;
        fc1_weights[44][146] = 16'sd-2;
        fc1_weights[44][147] = 16'sd79;
        fc1_weights[44][148] = 16'sd-1;
        fc1_weights[44][149] = 16'sd-18;
        fc1_weights[44][150] = 16'sd-86;
        fc1_weights[44][151] = 16'sd16;
        fc1_weights[44][152] = 16'sd-10;
        fc1_weights[44][153] = 16'sd26;
        fc1_weights[44][154] = 16'sd-29;
        fc1_weights[44][155] = 16'sd43;
        fc1_weights[44][156] = 16'sd13;
        fc1_weights[44][157] = 16'sd34;
        fc1_weights[44][158] = 16'sd11;
        fc1_weights[44][159] = 16'sd66;
        fc1_weights[44][160] = 16'sd-47;
        fc1_weights[44][161] = 16'sd25;
        fc1_weights[44][162] = 16'sd16;
        fc1_weights[44][163] = 16'sd-11;
        fc1_weights[44][164] = 16'sd15;
        fc1_weights[44][165] = 16'sd-64;
        fc1_weights[44][166] = 16'sd-24;
        fc1_weights[44][167] = 16'sd-12;
        fc1_weights[44][168] = 16'sd-57;
        fc1_weights[44][169] = 16'sd-14;
        fc1_weights[44][170] = 16'sd-30;
        fc1_weights[44][171] = 16'sd28;
        fc1_weights[44][172] = 16'sd-10;
        fc1_weights[44][173] = 16'sd26;
        fc1_weights[44][174] = 16'sd10;
        fc1_weights[44][175] = 16'sd36;
        fc1_weights[44][176] = 16'sd-1;
        fc1_weights[44][177] = 16'sd0;
        fc1_weights[44][178] = 16'sd4;
        fc1_weights[44][179] = 16'sd3;
        fc1_weights[44][180] = 16'sd-19;
        fc1_weights[44][181] = 16'sd0;
        fc1_weights[44][182] = 16'sd-4;
        fc1_weights[44][183] = 16'sd22;
        fc1_weights[44][184] = 16'sd13;
        fc1_weights[44][185] = 16'sd55;
        fc1_weights[44][186] = 16'sd9;
        fc1_weights[44][187] = 16'sd-30;
        fc1_weights[44][188] = 16'sd-22;
        fc1_weights[44][189] = 16'sd-8;
        fc1_weights[44][190] = 16'sd33;
        fc1_weights[44][191] = 16'sd-20;
        fc1_weights[44][192] = 16'sd-73;
        fc1_weights[44][193] = 16'sd-52;
        fc1_weights[44][194] = 16'sd-28;
        fc1_weights[44][195] = 16'sd-53;
        fc1_weights[44][196] = 16'sd-3;
        fc1_weights[44][197] = 16'sd-15;
        fc1_weights[44][198] = 16'sd-30;
        fc1_weights[44][199] = 16'sd17;
        fc1_weights[44][200] = 16'sd29;
        fc1_weights[44][201] = 16'sd-7;
        fc1_weights[44][202] = 16'sd24;
        fc1_weights[44][203] = 16'sd18;
        fc1_weights[44][204] = 16'sd-11;
        fc1_weights[44][205] = 16'sd20;
        fc1_weights[44][206] = 16'sd-38;
        fc1_weights[44][207] = 16'sd-17;
        fc1_weights[45][0] = 16'sd-26;
        fc1_weights[45][1] = 16'sd-16;
        fc1_weights[45][2] = 16'sd-83;
        fc1_weights[45][3] = 16'sd-19;
        fc1_weights[45][4] = 16'sd-7;
        fc1_weights[45][5] = 16'sd-25;
        fc1_weights[45][6] = 16'sd-49;
        fc1_weights[45][7] = 16'sd39;
        fc1_weights[45][8] = 16'sd-9;
        fc1_weights[45][9] = 16'sd-31;
        fc1_weights[45][10] = 16'sd18;
        fc1_weights[45][11] = 16'sd15;
        fc1_weights[45][12] = 16'sd1;
        fc1_weights[45][13] = 16'sd-64;
        fc1_weights[45][14] = 16'sd-85;
        fc1_weights[45][15] = 16'sd-23;
        fc1_weights[45][16] = 16'sd-140;
        fc1_weights[45][17] = 16'sd-107;
        fc1_weights[45][18] = 16'sd-56;
        fc1_weights[45][19] = 16'sd-52;
        fc1_weights[45][20] = 16'sd28;
        fc1_weights[45][21] = 16'sd-16;
        fc1_weights[45][22] = 16'sd-50;
        fc1_weights[45][23] = 16'sd-2;
        fc1_weights[45][24] = 16'sd10;
        fc1_weights[45][25] = 16'sd42;
        fc1_weights[45][26] = 16'sd-19;
        fc1_weights[45][27] = 16'sd-9;
        fc1_weights[45][28] = 16'sd26;
        fc1_weights[45][29] = 16'sd28;
        fc1_weights[45][30] = 16'sd-44;
        fc1_weights[45][31] = 16'sd43;
        fc1_weights[45][32] = 16'sd3;
        fc1_weights[45][33] = 16'sd13;
        fc1_weights[45][34] = 16'sd2;
        fc1_weights[45][35] = 16'sd-23;
        fc1_weights[45][36] = 16'sd53;
        fc1_weights[45][37] = 16'sd118;
        fc1_weights[45][38] = 16'sd12;
        fc1_weights[45][39] = 16'sd-78;
        fc1_weights[45][40] = 16'sd27;
        fc1_weights[45][41] = 16'sd-42;
        fc1_weights[45][42] = 16'sd-16;
        fc1_weights[45][43] = 16'sd-37;
        fc1_weights[45][44] = 16'sd3;
        fc1_weights[45][45] = 16'sd-22;
        fc1_weights[45][46] = 16'sd10;
        fc1_weights[45][47] = 16'sd32;
        fc1_weights[45][48] = 16'sd33;
        fc1_weights[45][49] = 16'sd57;
        fc1_weights[45][50] = 16'sd-6;
        fc1_weights[45][51] = 16'sd10;
        fc1_weights[45][52] = 16'sd11;
        fc1_weights[45][53] = 16'sd-11;
        fc1_weights[45][54] = 16'sd79;
        fc1_weights[45][55] = 16'sd-22;
        fc1_weights[45][56] = 16'sd-58;
        fc1_weights[45][57] = 16'sd-19;
        fc1_weights[45][58] = 16'sd-22;
        fc1_weights[45][59] = 16'sd21;
        fc1_weights[45][60] = 16'sd74;
        fc1_weights[45][61] = 16'sd42;
        fc1_weights[45][62] = 16'sd38;
        fc1_weights[45][63] = 16'sd16;
        fc1_weights[45][64] = 16'sd43;
        fc1_weights[45][65] = 16'sd-17;
        fc1_weights[45][66] = 16'sd-101;
        fc1_weights[45][67] = 16'sd-103;
        fc1_weights[45][68] = 16'sd-94;
        fc1_weights[45][69] = 16'sd-2;
        fc1_weights[45][70] = 16'sd-29;
        fc1_weights[45][71] = 16'sd20;
        fc1_weights[45][72] = 16'sd47;
        fc1_weights[45][73] = 16'sd-36;
        fc1_weights[45][74] = 16'sd18;
        fc1_weights[45][75] = 16'sd-54;
        fc1_weights[45][76] = 16'sd9;
        fc1_weights[45][77] = 16'sd7;
        fc1_weights[45][78] = 16'sd-1;
        fc1_weights[45][79] = 16'sd109;
        fc1_weights[45][80] = 16'sd-59;
        fc1_weights[45][81] = 16'sd-7;
        fc1_weights[45][82] = 16'sd-29;
        fc1_weights[45][83] = 16'sd7;
        fc1_weights[45][84] = 16'sd1;
        fc1_weights[45][85] = 16'sd-86;
        fc1_weights[45][86] = 16'sd23;
        fc1_weights[45][87] = 16'sd32;
        fc1_weights[45][88] = 16'sd34;
        fc1_weights[45][89] = 16'sd28;
        fc1_weights[45][90] = 16'sd37;
        fc1_weights[45][91] = 16'sd-28;
        fc1_weights[45][92] = 16'sd84;
        fc1_weights[45][93] = 16'sd-80;
        fc1_weights[45][94] = 16'sd-129;
        fc1_weights[45][95] = 16'sd-73;
        fc1_weights[45][96] = 16'sd-56;
        fc1_weights[45][97] = 16'sd4;
        fc1_weights[45][98] = 16'sd-34;
        fc1_weights[45][99] = 16'sd-45;
        fc1_weights[45][100] = 16'sd15;
        fc1_weights[45][101] = 16'sd-3;
        fc1_weights[45][102] = 16'sd-81;
        fc1_weights[45][103] = 16'sd-138;
        fc1_weights[45][104] = 16'sd138;
        fc1_weights[45][105] = 16'sd4;
        fc1_weights[45][106] = 16'sd72;
        fc1_weights[45][107] = 16'sd20;
        fc1_weights[45][108] = 16'sd-15;
        fc1_weights[45][109] = 16'sd-72;
        fc1_weights[45][110] = 16'sd-57;
        fc1_weights[45][111] = 16'sd-19;
        fc1_weights[45][112] = 16'sd61;
        fc1_weights[45][113] = 16'sd97;
        fc1_weights[45][114] = 16'sd41;
        fc1_weights[45][115] = 16'sd27;
        fc1_weights[45][116] = 16'sd120;
        fc1_weights[45][117] = 16'sd61;
        fc1_weights[45][118] = 16'sd9;
        fc1_weights[45][119] = 16'sd45;
        fc1_weights[45][120] = 16'sd-24;
        fc1_weights[45][121] = 16'sd39;
        fc1_weights[45][122] = 16'sd-9;
        fc1_weights[45][123] = 16'sd49;
        fc1_weights[45][124] = 16'sd-42;
        fc1_weights[45][125] = 16'sd5;
        fc1_weights[45][126] = 16'sd-40;
        fc1_weights[45][127] = 16'sd0;
        fc1_weights[45][128] = 16'sd19;
        fc1_weights[45][129] = 16'sd-31;
        fc1_weights[45][130] = 16'sd34;
        fc1_weights[45][131] = 16'sd-46;
        fc1_weights[45][132] = 16'sd-36;
        fc1_weights[45][133] = 16'sd-100;
        fc1_weights[45][134] = 16'sd-52;
        fc1_weights[45][135] = 16'sd-65;
        fc1_weights[45][136] = 16'sd-12;
        fc1_weights[45][137] = 16'sd39;
        fc1_weights[45][138] = 16'sd51;
        fc1_weights[45][139] = 16'sd54;
        fc1_weights[45][140] = 16'sd27;
        fc1_weights[45][141] = 16'sd-41;
        fc1_weights[45][142] = 16'sd0;
        fc1_weights[45][143] = 16'sd-36;
        fc1_weights[45][144] = 16'sd-49;
        fc1_weights[45][145] = 16'sd35;
        fc1_weights[45][146] = 16'sd44;
        fc1_weights[45][147] = 16'sd18;
        fc1_weights[45][148] = 16'sd68;
        fc1_weights[45][149] = 16'sd1;
        fc1_weights[45][150] = 16'sd-11;
        fc1_weights[45][151] = 16'sd36;
        fc1_weights[45][152] = 16'sd14;
        fc1_weights[45][153] = 16'sd63;
        fc1_weights[45][154] = 16'sd-65;
        fc1_weights[45][155] = 16'sd-2;
        fc1_weights[45][156] = 16'sd39;
        fc1_weights[45][157] = 16'sd43;
        fc1_weights[45][158] = 16'sd-21;
        fc1_weights[45][159] = 16'sd88;
        fc1_weights[45][160] = 16'sd-60;
        fc1_weights[45][161] = 16'sd-38;
        fc1_weights[45][162] = 16'sd22;
        fc1_weights[45][163] = 16'sd-16;
        fc1_weights[45][164] = 16'sd42;
        fc1_weights[45][165] = 16'sd-85;
        fc1_weights[45][166] = 16'sd27;
        fc1_weights[45][167] = 16'sd-54;
        fc1_weights[45][168] = 16'sd53;
        fc1_weights[45][169] = 16'sd-56;
        fc1_weights[45][170] = 16'sd-42;
        fc1_weights[45][171] = 16'sd17;
        fc1_weights[45][172] = 16'sd28;
        fc1_weights[45][173] = 16'sd21;
        fc1_weights[45][174] = 16'sd12;
        fc1_weights[45][175] = 16'sd46;
        fc1_weights[45][176] = 16'sd-4;
        fc1_weights[45][177] = 16'sd60;
        fc1_weights[45][178] = 16'sd-37;
        fc1_weights[45][179] = 16'sd-7;
        fc1_weights[45][180] = 16'sd19;
        fc1_weights[45][181] = 16'sd58;
        fc1_weights[45][182] = 16'sd7;
        fc1_weights[45][183] = 16'sd-19;
        fc1_weights[45][184] = 16'sd-13;
        fc1_weights[45][185] = 16'sd118;
        fc1_weights[45][186] = 16'sd-11;
        fc1_weights[45][187] = 16'sd13;
        fc1_weights[45][188] = 16'sd18;
        fc1_weights[45][189] = 16'sd70;
        fc1_weights[45][190] = 16'sd56;
        fc1_weights[45][191] = 16'sd14;
        fc1_weights[45][192] = 16'sd-106;
        fc1_weights[45][193] = 16'sd-71;
        fc1_weights[45][194] = 16'sd-26;
        fc1_weights[45][195] = 16'sd33;
        fc1_weights[45][196] = 16'sd-18;
        fc1_weights[45][197] = 16'sd32;
        fc1_weights[45][198] = 16'sd-71;
        fc1_weights[45][199] = 16'sd52;
        fc1_weights[45][200] = 16'sd40;
        fc1_weights[45][201] = 16'sd37;
        fc1_weights[45][202] = 16'sd-3;
        fc1_weights[45][203] = 16'sd49;
        fc1_weights[45][204] = 16'sd47;
        fc1_weights[45][205] = 16'sd81;
        fc1_weights[45][206] = 16'sd18;
        fc1_weights[45][207] = 16'sd-9;
        fc1_weights[46][0] = 16'sd40;
        fc1_weights[46][1] = 16'sd23;
        fc1_weights[46][2] = 16'sd20;
        fc1_weights[46][3] = 16'sd-38;
        fc1_weights[46][4] = 16'sd-34;
        fc1_weights[46][5] = 16'sd17;
        fc1_weights[46][6] = 16'sd15;
        fc1_weights[46][7] = 16'sd38;
        fc1_weights[46][8] = 16'sd-62;
        fc1_weights[46][9] = 16'sd-65;
        fc1_weights[46][10] = 16'sd-58;
        fc1_weights[46][11] = 16'sd-120;
        fc1_weights[46][12] = 16'sd-76;
        fc1_weights[46][13] = 16'sd8;
        fc1_weights[46][14] = 16'sd96;
        fc1_weights[46][15] = 16'sd134;
        fc1_weights[46][16] = 16'sd77;
        fc1_weights[46][17] = 16'sd15;
        fc1_weights[46][18] = 16'sd46;
        fc1_weights[46][19] = 16'sd38;
        fc1_weights[46][20] = 16'sd29;
        fc1_weights[46][21] = 16'sd-5;
        fc1_weights[46][22] = 16'sd-15;
        fc1_weights[46][23] = 16'sd22;
        fc1_weights[46][24] = 16'sd-33;
        fc1_weights[46][25] = 16'sd20;
        fc1_weights[46][26] = 16'sd21;
        fc1_weights[46][27] = 16'sd19;
        fc1_weights[46][28] = 16'sd1;
        fc1_weights[46][29] = 16'sd21;
        fc1_weights[46][30] = 16'sd14;
        fc1_weights[46][31] = 16'sd3;
        fc1_weights[46][32] = 16'sd-10;
        fc1_weights[46][33] = 16'sd-46;
        fc1_weights[46][34] = 16'sd-50;
        fc1_weights[46][35] = 16'sd-62;
        fc1_weights[46][36] = 16'sd-19;
        fc1_weights[46][37] = 16'sd-64;
        fc1_weights[46][38] = 16'sd-11;
        fc1_weights[46][39] = 16'sd-31;
        fc1_weights[46][40] = 16'sd110;
        fc1_weights[46][41] = 16'sd106;
        fc1_weights[46][42] = 16'sd-41;
        fc1_weights[46][43] = 16'sd-26;
        fc1_weights[46][44] = 16'sd-12;
        fc1_weights[46][45] = 16'sd-117;
        fc1_weights[46][46] = 16'sd-23;
        fc1_weights[46][47] = 16'sd-56;
        fc1_weights[46][48] = 16'sd-19;
        fc1_weights[46][49] = 16'sd20;
        fc1_weights[46][50] = 16'sd19;
        fc1_weights[46][51] = 16'sd-33;
        fc1_weights[46][52] = 16'sd25;
        fc1_weights[46][53] = 16'sd21;
        fc1_weights[46][54] = 16'sd2;
        fc1_weights[46][55] = 16'sd63;
        fc1_weights[46][56] = 16'sd41;
        fc1_weights[46][57] = 16'sd30;
        fc1_weights[46][58] = 16'sd49;
        fc1_weights[46][59] = 16'sd10;
        fc1_weights[46][60] = 16'sd26;
        fc1_weights[46][61] = 16'sd-26;
        fc1_weights[46][62] = 16'sd-55;
        fc1_weights[46][63] = 16'sd13;
        fc1_weights[46][64] = 16'sd18;
        fc1_weights[46][65] = 16'sd-39;
        fc1_weights[46][66] = 16'sd53;
        fc1_weights[46][67] = 16'sd41;
        fc1_weights[46][68] = 16'sd10;
        fc1_weights[46][69] = 16'sd-13;
        fc1_weights[46][70] = 16'sd55;
        fc1_weights[46][71] = 16'sd24;
        fc1_weights[46][72] = 16'sd-6;
        fc1_weights[46][73] = 16'sd5;
        fc1_weights[46][74] = 16'sd-13;
        fc1_weights[46][75] = 16'sd-20;
        fc1_weights[46][76] = 16'sd-9;
        fc1_weights[46][77] = 16'sd-23;
        fc1_weights[46][78] = 16'sd-28;
        fc1_weights[46][79] = 16'sd24;
        fc1_weights[46][80] = 16'sd-4;
        fc1_weights[46][81] = 16'sd31;
        fc1_weights[46][82] = 16'sd-63;
        fc1_weights[46][83] = 16'sd40;
        fc1_weights[46][84] = 16'sd16;
        fc1_weights[46][85] = 16'sd-21;
        fc1_weights[46][86] = 16'sd-71;
        fc1_weights[46][87] = 16'sd-32;
        fc1_weights[46][88] = 16'sd-62;
        fc1_weights[46][89] = 16'sd-3;
        fc1_weights[46][90] = 16'sd43;
        fc1_weights[46][91] = 16'sd31;
        fc1_weights[46][92] = 16'sd52;
        fc1_weights[46][93] = 16'sd105;
        fc1_weights[46][94] = 16'sd-27;
        fc1_weights[46][95] = 16'sd-47;
        fc1_weights[46][96] = 16'sd-4;
        fc1_weights[46][97] = 16'sd27;
        fc1_weights[46][98] = 16'sd54;
        fc1_weights[46][99] = 16'sd-9;
        fc1_weights[46][100] = 16'sd17;
        fc1_weights[46][101] = 16'sd2;
        fc1_weights[46][102] = 16'sd-31;
        fc1_weights[46][103] = 16'sd-24;
        fc1_weights[46][104] = 16'sd48;
        fc1_weights[46][105] = 16'sd-34;
        fc1_weights[46][106] = 16'sd28;
        fc1_weights[46][107] = 16'sd-26;
        fc1_weights[46][108] = 16'sd8;
        fc1_weights[46][109] = 16'sd51;
        fc1_weights[46][110] = 16'sd44;
        fc1_weights[46][111] = 16'sd-56;
        fc1_weights[46][112] = 16'sd-20;
        fc1_weights[46][113] = 16'sd-10;
        fc1_weights[46][114] = 16'sd-1;
        fc1_weights[46][115] = 16'sd-66;
        fc1_weights[46][116] = 16'sd-37;
        fc1_weights[46][117] = 16'sd-26;
        fc1_weights[46][118] = 16'sd-11;
        fc1_weights[46][119] = 16'sd-12;
        fc1_weights[46][120] = 16'sd-16;
        fc1_weights[46][121] = 16'sd-25;
        fc1_weights[46][122] = 16'sd-75;
        fc1_weights[46][123] = 16'sd-61;
        fc1_weights[46][124] = 16'sd-60;
        fc1_weights[46][125] = 16'sd-98;
        fc1_weights[46][126] = 16'sd-88;
        fc1_weights[46][127] = 16'sd-15;
        fc1_weights[46][128] = 16'sd-37;
        fc1_weights[46][129] = 16'sd-46;
        fc1_weights[46][130] = 16'sd-44;
        fc1_weights[46][131] = 16'sd13;
        fc1_weights[46][132] = 16'sd-7;
        fc1_weights[46][133] = 16'sd70;
        fc1_weights[46][134] = 16'sd42;
        fc1_weights[46][135] = 16'sd58;
        fc1_weights[46][136] = 16'sd108;
        fc1_weights[46][137] = 16'sd3;
        fc1_weights[46][138] = 16'sd74;
        fc1_weights[46][139] = 16'sd-83;
        fc1_weights[46][140] = 16'sd-62;
        fc1_weights[46][141] = 16'sd7;
        fc1_weights[46][142] = 16'sd-40;
        fc1_weights[46][143] = 16'sd-29;
        fc1_weights[46][144] = 16'sd64;
        fc1_weights[46][145] = 16'sd-17;
        fc1_weights[46][146] = 16'sd47;
        fc1_weights[46][147] = 16'sd103;
        fc1_weights[46][148] = 16'sd13;
        fc1_weights[46][149] = 16'sd-29;
        fc1_weights[46][150] = 16'sd2;
        fc1_weights[46][151] = 16'sd-12;
        fc1_weights[46][152] = 16'sd-10;
        fc1_weights[46][153] = 16'sd-13;
        fc1_weights[46][154] = 16'sd20;
        fc1_weights[46][155] = 16'sd28;
        fc1_weights[46][156] = 16'sd36;
        fc1_weights[46][157] = 16'sd63;
        fc1_weights[46][158] = 16'sd32;
        fc1_weights[46][159] = 16'sd57;
        fc1_weights[46][160] = 16'sd27;
        fc1_weights[46][161] = 16'sd16;
        fc1_weights[46][162] = 16'sd21;
        fc1_weights[46][163] = 16'sd18;
        fc1_weights[46][164] = 16'sd-54;
        fc1_weights[46][165] = 16'sd10;
        fc1_weights[46][166] = 16'sd-11;
        fc1_weights[46][167] = 16'sd15;
        fc1_weights[46][168] = 16'sd-7;
        fc1_weights[46][169] = 16'sd4;
        fc1_weights[46][170] = 16'sd14;
        fc1_weights[46][171] = 16'sd-39;
        fc1_weights[46][172] = 16'sd24;
        fc1_weights[46][173] = 16'sd-28;
        fc1_weights[46][174] = 16'sd1;
        fc1_weights[46][175] = 16'sd10;
        fc1_weights[46][176] = 16'sd20;
        fc1_weights[46][177] = 16'sd-35;
        fc1_weights[46][178] = 16'sd12;
        fc1_weights[46][179] = 16'sd20;
        fc1_weights[46][180] = 16'sd15;
        fc1_weights[46][181] = 16'sd48;
        fc1_weights[46][182] = 16'sd2;
        fc1_weights[46][183] = 16'sd66;
        fc1_weights[46][184] = 16'sd18;
        fc1_weights[46][185] = 16'sd-9;
        fc1_weights[46][186] = 16'sd-10;
        fc1_weights[46][187] = 16'sd-25;
        fc1_weights[46][188] = 16'sd-79;
        fc1_weights[46][189] = 16'sd-54;
        fc1_weights[46][190] = 16'sd40;
        fc1_weights[46][191] = 16'sd-3;
        fc1_weights[46][192] = 16'sd-12;
        fc1_weights[46][193] = 16'sd-11;
        fc1_weights[46][194] = 16'sd3;
        fc1_weights[46][195] = 16'sd16;
        fc1_weights[46][196] = 16'sd-13;
        fc1_weights[46][197] = 16'sd8;
        fc1_weights[46][198] = 16'sd-46;
        fc1_weights[46][199] = 16'sd-20;
        fc1_weights[46][200] = 16'sd-7;
        fc1_weights[46][201] = 16'sd-61;
        fc1_weights[46][202] = 16'sd-46;
        fc1_weights[46][203] = 16'sd23;
        fc1_weights[46][204] = 16'sd6;
        fc1_weights[46][205] = 16'sd48;
        fc1_weights[46][206] = 16'sd-21;
        fc1_weights[46][207] = 16'sd67;
        fc1_weights[47][0] = 16'sd20;
        fc1_weights[47][1] = 16'sd13;
        fc1_weights[47][2] = 16'sd-2;
        fc1_weights[47][3] = 16'sd-3;
        fc1_weights[47][4] = 16'sd-4;
        fc1_weights[47][5] = 16'sd-27;
        fc1_weights[47][6] = 16'sd-15;
        fc1_weights[47][7] = 16'sd-31;
        fc1_weights[47][8] = 16'sd19;
        fc1_weights[47][9] = 16'sd-8;
        fc1_weights[47][10] = 16'sd-37;
        fc1_weights[47][11] = 16'sd33;
        fc1_weights[47][12] = 16'sd38;
        fc1_weights[47][13] = 16'sd16;
        fc1_weights[47][14] = 16'sd-14;
        fc1_weights[47][15] = 16'sd-58;
        fc1_weights[47][16] = 16'sd5;
        fc1_weights[47][17] = 16'sd-9;
        fc1_weights[47][18] = 16'sd-30;
        fc1_weights[47][19] = 16'sd12;
        fc1_weights[47][20] = 16'sd-27;
        fc1_weights[47][21] = 16'sd-14;
        fc1_weights[47][22] = 16'sd-13;
        fc1_weights[47][23] = 16'sd-13;
        fc1_weights[47][24] = 16'sd-30;
        fc1_weights[47][25] = 16'sd-46;
        fc1_weights[47][26] = 16'sd6;
        fc1_weights[47][27] = 16'sd15;
        fc1_weights[47][28] = 16'sd11;
        fc1_weights[47][29] = 16'sd-9;
        fc1_weights[47][30] = 16'sd-20;
        fc1_weights[47][31] = 16'sd-13;
        fc1_weights[47][32] = 16'sd0;
        fc1_weights[47][33] = 16'sd-5;
        fc1_weights[47][34] = 16'sd1;
        fc1_weights[47][35] = 16'sd-14;
        fc1_weights[47][36] = 16'sd-59;
        fc1_weights[47][37] = 16'sd-54;
        fc1_weights[47][38] = 16'sd-14;
        fc1_weights[47][39] = 16'sd26;
        fc1_weights[47][40] = 16'sd-25;
        fc1_weights[47][41] = 16'sd-10;
        fc1_weights[47][42] = 16'sd8;
        fc1_weights[47][43] = 16'sd26;
        fc1_weights[47][44] = 16'sd-26;
        fc1_weights[47][45] = 16'sd-2;
        fc1_weights[47][46] = 16'sd8;
        fc1_weights[47][47] = 16'sd21;
        fc1_weights[47][48] = 16'sd-42;
        fc1_weights[47][49] = 16'sd-43;
        fc1_weights[47][50] = 16'sd-20;
        fc1_weights[47][51] = 16'sd26;
        fc1_weights[47][52] = 16'sd-5;
        fc1_weights[47][53] = 16'sd-9;
        fc1_weights[47][54] = 16'sd-8;
        fc1_weights[47][55] = 16'sd-19;
        fc1_weights[47][56] = 16'sd-34;
        fc1_weights[47][57] = 16'sd-44;
        fc1_weights[47][58] = 16'sd-2;
        fc1_weights[47][59] = 16'sd-6;
        fc1_weights[47][60] = 16'sd-26;
        fc1_weights[47][61] = 16'sd-1;
        fc1_weights[47][62] = 16'sd5;
        fc1_weights[47][63] = 16'sd-54;
        fc1_weights[47][64] = 16'sd-3;
        fc1_weights[47][65] = 16'sd60;
        fc1_weights[47][66] = 16'sd-13;
        fc1_weights[47][67] = 16'sd3;
        fc1_weights[47][68] = 16'sd-10;
        fc1_weights[47][69] = 16'sd-24;
        fc1_weights[47][70] = 16'sd-43;
        fc1_weights[47][71] = 16'sd12;
        fc1_weights[47][72] = 16'sd-5;
        fc1_weights[47][73] = 16'sd-21;
        fc1_weights[47][74] = 16'sd-13;
        fc1_weights[47][75] = 16'sd-5;
        fc1_weights[47][76] = 16'sd-9;
        fc1_weights[47][77] = 16'sd-5;
        fc1_weights[47][78] = 16'sd4;
        fc1_weights[47][79] = 16'sd0;
        fc1_weights[47][80] = 16'sd2;
        fc1_weights[47][81] = 16'sd-11;
        fc1_weights[47][82] = 16'sd-2;
        fc1_weights[47][83] = 16'sd-14;
        fc1_weights[47][84] = 16'sd-15;
        fc1_weights[47][85] = 16'sd6;
        fc1_weights[47][86] = 16'sd-21;
        fc1_weights[47][87] = 16'sd-22;
        fc1_weights[47][88] = 16'sd6;
        fc1_weights[47][89] = 16'sd-2;
        fc1_weights[47][90] = 16'sd43;
        fc1_weights[47][91] = 16'sd-2;
        fc1_weights[47][92] = 16'sd9;
        fc1_weights[47][93] = 16'sd-36;
        fc1_weights[47][94] = 16'sd-1;
        fc1_weights[47][95] = 16'sd7;
        fc1_weights[47][96] = 16'sd4;
        fc1_weights[47][97] = 16'sd21;
        fc1_weights[47][98] = 16'sd9;
        fc1_weights[47][99] = 16'sd16;
        fc1_weights[47][100] = 16'sd-1;
        fc1_weights[47][101] = 16'sd-25;
        fc1_weights[47][102] = 16'sd34;
        fc1_weights[47][103] = 16'sd35;
        fc1_weights[47][104] = 16'sd-22;
        fc1_weights[47][105] = 16'sd9;
        fc1_weights[47][106] = 16'sd-7;
        fc1_weights[47][107] = 16'sd-1;
        fc1_weights[47][108] = 16'sd-8;
        fc1_weights[47][109] = 16'sd-22;
        fc1_weights[47][110] = 16'sd-28;
        fc1_weights[47][111] = 16'sd-18;
        fc1_weights[47][112] = 16'sd-19;
        fc1_weights[47][113] = 16'sd27;
        fc1_weights[47][114] = 16'sd-43;
        fc1_weights[47][115] = 16'sd-28;
        fc1_weights[47][116] = 16'sd3;
        fc1_weights[47][117] = 16'sd7;
        fc1_weights[47][118] = 16'sd-18;
        fc1_weights[47][119] = 16'sd20;
        fc1_weights[47][120] = 16'sd34;
        fc1_weights[47][121] = 16'sd8;
        fc1_weights[47][122] = 16'sd19;
        fc1_weights[47][123] = 16'sd12;
        fc1_weights[47][124] = 16'sd14;
        fc1_weights[47][125] = 16'sd24;
        fc1_weights[47][126] = 16'sd10;
        fc1_weights[47][127] = 16'sd20;
        fc1_weights[47][128] = 16'sd-14;
        fc1_weights[47][129] = 16'sd19;
        fc1_weights[47][130] = 16'sd-37;
        fc1_weights[47][131] = 16'sd-11;
        fc1_weights[47][132] = 16'sd-4;
        fc1_weights[47][133] = 16'sd10;
        fc1_weights[47][134] = 16'sd34;
        fc1_weights[47][135] = 16'sd5;
        fc1_weights[47][136] = 16'sd-17;
        fc1_weights[47][137] = 16'sd-10;
        fc1_weights[47][138] = 16'sd-11;
        fc1_weights[47][139] = 16'sd11;
        fc1_weights[47][140] = 16'sd4;
        fc1_weights[47][141] = 16'sd-6;
        fc1_weights[47][142] = 16'sd10;
        fc1_weights[47][143] = 16'sd-32;
        fc1_weights[47][144] = 16'sd5;
        fc1_weights[47][145] = 16'sd3;
        fc1_weights[47][146] = 16'sd-14;
        fc1_weights[47][147] = 16'sd-24;
        fc1_weights[47][148] = 16'sd8;
        fc1_weights[47][149] = 16'sd28;
        fc1_weights[47][150] = 16'sd30;
        fc1_weights[47][151] = 16'sd46;
        fc1_weights[47][152] = 16'sd55;
        fc1_weights[47][153] = 16'sd25;
        fc1_weights[47][154] = 16'sd32;
        fc1_weights[47][155] = 16'sd23;
        fc1_weights[47][156] = 16'sd16;
        fc1_weights[47][157] = 16'sd6;
        fc1_weights[47][158] = 16'sd28;
        fc1_weights[47][159] = 16'sd15;
        fc1_weights[47][160] = 16'sd-12;
        fc1_weights[47][161] = 16'sd20;
        fc1_weights[47][162] = 16'sd-5;
        fc1_weights[47][163] = 16'sd4;
        fc1_weights[47][164] = 16'sd2;
        fc1_weights[47][165] = 16'sd27;
        fc1_weights[47][166] = 16'sd-7;
        fc1_weights[47][167] = 16'sd12;
        fc1_weights[47][168] = 16'sd-15;
        fc1_weights[47][169] = 16'sd9;
        fc1_weights[47][170] = 16'sd6;
        fc1_weights[47][171] = 16'sd16;
        fc1_weights[47][172] = 16'sd12;
        fc1_weights[47][173] = 16'sd43;
        fc1_weights[47][174] = 16'sd28;
        fc1_weights[47][175] = 16'sd34;
        fc1_weights[47][176] = 16'sd29;
        fc1_weights[47][177] = 16'sd45;
        fc1_weights[47][178] = 16'sd47;
        fc1_weights[47][179] = 16'sd39;
        fc1_weights[47][180] = 16'sd48;
        fc1_weights[47][181] = 16'sd15;
        fc1_weights[47][182] = 16'sd-8;
        fc1_weights[47][183] = 16'sd-9;
        fc1_weights[47][184] = 16'sd-1;
        fc1_weights[47][185] = 16'sd-23;
        fc1_weights[47][186] = 16'sd-7;
        fc1_weights[47][187] = 16'sd-8;
        fc1_weights[47][188] = 16'sd-5;
        fc1_weights[47][189] = 16'sd-22;
        fc1_weights[47][190] = 16'sd27;
        fc1_weights[47][191] = 16'sd-11;
        fc1_weights[47][192] = 16'sd11;
        fc1_weights[47][193] = 16'sd5;
        fc1_weights[47][194] = 16'sd23;
        fc1_weights[47][195] = 16'sd11;
        fc1_weights[47][196] = 16'sd6;
        fc1_weights[47][197] = 16'sd28;
        fc1_weights[47][198] = 16'sd34;
        fc1_weights[47][199] = 16'sd34;
        fc1_weights[47][200] = 16'sd15;
        fc1_weights[47][201] = 16'sd19;
        fc1_weights[47][202] = 16'sd31;
        fc1_weights[47][203] = 16'sd13;
        fc1_weights[47][204] = 16'sd27;
        fc1_weights[47][205] = 16'sd3;
        fc1_weights[47][206] = 16'sd32;
        fc1_weights[47][207] = 16'sd4;
        fc1_weights[48][0] = 16'sd-2;
        fc1_weights[48][1] = 16'sd10;
        fc1_weights[48][2] = 16'sd24;
        fc1_weights[48][3] = 16'sd7;
        fc1_weights[48][4] = 16'sd1;
        fc1_weights[48][5] = 16'sd-9;
        fc1_weights[48][6] = 16'sd-20;
        fc1_weights[48][7] = 16'sd24;
        fc1_weights[48][8] = 16'sd2;
        fc1_weights[48][9] = 16'sd-10;
        fc1_weights[48][10] = 16'sd-37;
        fc1_weights[48][11] = 16'sd-27;
        fc1_weights[48][12] = 16'sd-40;
        fc1_weights[48][13] = 16'sd-41;
        fc1_weights[48][14] = 16'sd7;
        fc1_weights[48][15] = 16'sd24;
        fc1_weights[48][16] = 16'sd-10;
        fc1_weights[48][17] = 16'sd26;
        fc1_weights[48][18] = 16'sd-3;
        fc1_weights[48][19] = 16'sd-5;
        fc1_weights[48][20] = 16'sd1;
        fc1_weights[48][21] = 16'sd-8;
        fc1_weights[48][22] = 16'sd15;
        fc1_weights[48][23] = 16'sd32;
        fc1_weights[48][24] = 16'sd32;
        fc1_weights[48][25] = 16'sd49;
        fc1_weights[48][26] = 16'sd12;
        fc1_weights[48][27] = 16'sd5;
        fc1_weights[48][28] = 16'sd11;
        fc1_weights[48][29] = 16'sd35;
        fc1_weights[48][30] = 16'sd18;
        fc1_weights[48][31] = 16'sd50;
        fc1_weights[48][32] = 16'sd14;
        fc1_weights[48][33] = 16'sd17;
        fc1_weights[48][34] = 16'sd10;
        fc1_weights[48][35] = 16'sd-1;
        fc1_weights[48][36] = 16'sd-22;
        fc1_weights[48][37] = 16'sd24;
        fc1_weights[48][38] = 16'sd-14;
        fc1_weights[48][39] = 16'sd14;
        fc1_weights[48][40] = 16'sd-6;
        fc1_weights[48][41] = 16'sd-17;
        fc1_weights[48][42] = 16'sd19;
        fc1_weights[48][43] = 16'sd-34;
        fc1_weights[48][44] = 16'sd-41;
        fc1_weights[48][45] = 16'sd-74;
        fc1_weights[48][46] = 16'sd-34;
        fc1_weights[48][47] = 16'sd-9;
        fc1_weights[48][48] = 16'sd-13;
        fc1_weights[48][49] = 16'sd1;
        fc1_weights[48][50] = 16'sd17;
        fc1_weights[48][51] = 16'sd-20;
        fc1_weights[48][52] = 16'sd31;
        fc1_weights[48][53] = 16'sd59;
        fc1_weights[48][54] = 16'sd-16;
        fc1_weights[48][55] = 16'sd-2;
        fc1_weights[48][56] = 16'sd1;
        fc1_weights[48][57] = 16'sd20;
        fc1_weights[48][58] = 16'sd4;
        fc1_weights[48][59] = 16'sd37;
        fc1_weights[48][60] = 16'sd3;
        fc1_weights[48][61] = 16'sd24;
        fc1_weights[48][62] = 16'sd-50;
        fc1_weights[48][63] = 16'sd-12;
        fc1_weights[48][64] = 16'sd8;
        fc1_weights[48][65] = 16'sd-44;
        fc1_weights[48][66] = 16'sd-29;
        fc1_weights[48][67] = 16'sd11;
        fc1_weights[48][68] = 16'sd31;
        fc1_weights[48][69] = 16'sd3;
        fc1_weights[48][70] = 16'sd-14;
        fc1_weights[48][71] = 16'sd-24;
        fc1_weights[48][72] = 16'sd-32;
        fc1_weights[48][73] = 16'sd6;
        fc1_weights[48][74] = 16'sd-2;
        fc1_weights[48][75] = 16'sd17;
        fc1_weights[48][76] = 16'sd19;
        fc1_weights[48][77] = 16'sd18;
        fc1_weights[48][78] = 16'sd33;
        fc1_weights[48][79] = 16'sd18;
        fc1_weights[48][80] = 16'sd5;
        fc1_weights[48][81] = 16'sd2;
        fc1_weights[48][82] = 16'sd26;
        fc1_weights[48][83] = 16'sd-8;
        fc1_weights[48][84] = 16'sd12;
        fc1_weights[48][85] = 16'sd19;
        fc1_weights[48][86] = 16'sd27;
        fc1_weights[48][87] = 16'sd3;
        fc1_weights[48][88] = 16'sd-62;
        fc1_weights[48][89] = 16'sd-40;
        fc1_weights[48][90] = 16'sd-14;
        fc1_weights[48][91] = 16'sd-59;
        fc1_weights[48][92] = 16'sd-17;
        fc1_weights[48][93] = 16'sd13;
        fc1_weights[48][94] = 16'sd1;
        fc1_weights[48][95] = 16'sd-15;
        fc1_weights[48][96] = 16'sd-22;
        fc1_weights[48][97] = 16'sd20;
        fc1_weights[48][98] = 16'sd7;
        fc1_weights[48][99] = 16'sd9;
        fc1_weights[48][100] = 16'sd35;
        fc1_weights[48][101] = 16'sd37;
        fc1_weights[48][102] = 16'sd-2;
        fc1_weights[48][103] = 16'sd-18;
        fc1_weights[48][104] = 16'sd24;
        fc1_weights[48][105] = 16'sd-1;
        fc1_weights[48][106] = 16'sd1;
        fc1_weights[48][107] = 16'sd-36;
        fc1_weights[48][108] = 16'sd-32;
        fc1_weights[48][109] = 16'sd-17;
        fc1_weights[48][110] = 16'sd-9;
        fc1_weights[48][111] = 16'sd-10;
        fc1_weights[48][112] = 16'sd-24;
        fc1_weights[48][113] = 16'sd5;
        fc1_weights[48][114] = 16'sd-26;
        fc1_weights[48][115] = 16'sd19;
        fc1_weights[48][116] = 16'sd-29;
        fc1_weights[48][117] = 16'sd-53;
        fc1_weights[48][118] = 16'sd-21;
        fc1_weights[48][119] = 16'sd-26;
        fc1_weights[48][120] = 16'sd-64;
        fc1_weights[48][121] = 16'sd-4;
        fc1_weights[48][122] = 16'sd-61;
        fc1_weights[48][123] = 16'sd-20;
        fc1_weights[48][124] = 16'sd-16;
        fc1_weights[48][125] = 16'sd-36;
        fc1_weights[48][126] = 16'sd-23;
        fc1_weights[48][127] = 16'sd2;
        fc1_weights[48][128] = 16'sd-17;
        fc1_weights[48][129] = 16'sd-80;
        fc1_weights[48][130] = 16'sd-21;
        fc1_weights[48][131] = 16'sd-30;
        fc1_weights[48][132] = 16'sd-57;
        fc1_weights[48][133] = 16'sd-34;
        fc1_weights[48][134] = 16'sd-20;
        fc1_weights[48][135] = 16'sd-58;
        fc1_weights[48][136] = 16'sd-17;
        fc1_weights[48][137] = 16'sd-8;
        fc1_weights[48][138] = 16'sd11;
        fc1_weights[48][139] = 16'sd27;
        fc1_weights[48][140] = 16'sd-2;
        fc1_weights[48][141] = 16'sd50;
        fc1_weights[48][142] = 16'sd22;
        fc1_weights[48][143] = 16'sd2;
        fc1_weights[48][144] = 16'sd7;
        fc1_weights[48][145] = 16'sd2;
        fc1_weights[48][146] = 16'sd8;
        fc1_weights[48][147] = 16'sd39;
        fc1_weights[48][148] = 16'sd25;
        fc1_weights[48][149] = 16'sd-8;
        fc1_weights[48][150] = 16'sd9;
        fc1_weights[48][151] = 16'sd1;
        fc1_weights[48][152] = 16'sd21;
        fc1_weights[48][153] = 16'sd11;
        fc1_weights[48][154] = 16'sd-24;
        fc1_weights[48][155] = 16'sd3;
        fc1_weights[48][156] = 16'sd-12;
        fc1_weights[48][157] = 16'sd-22;
        fc1_weights[48][158] = 16'sd-23;
        fc1_weights[48][159] = 16'sd-61;
        fc1_weights[48][160] = 16'sd7;
        fc1_weights[48][161] = 16'sd38;
        fc1_weights[48][162] = 16'sd11;
        fc1_weights[48][163] = 16'sd-34;
        fc1_weights[48][164] = 16'sd-9;
        fc1_weights[48][165] = 16'sd-44;
        fc1_weights[48][166] = 16'sd4;
        fc1_weights[48][167] = 16'sd12;
        fc1_weights[48][168] = 16'sd23;
        fc1_weights[48][169] = 16'sd34;
        fc1_weights[48][170] = 16'sd47;
        fc1_weights[48][171] = 16'sd28;
        fc1_weights[48][172] = 16'sd18;
        fc1_weights[48][173] = 16'sd57;
        fc1_weights[48][174] = 16'sd36;
        fc1_weights[48][175] = 16'sd42;
        fc1_weights[48][176] = 16'sd19;
        fc1_weights[48][177] = 16'sd31;
        fc1_weights[48][178] = 16'sd8;
        fc1_weights[48][179] = 16'sd1;
        fc1_weights[48][180] = 16'sd-10;
        fc1_weights[48][181] = 16'sd-9;
        fc1_weights[48][182] = 16'sd11;
        fc1_weights[48][183] = 16'sd-8;
        fc1_weights[48][184] = 16'sd-48;
        fc1_weights[48][185] = 16'sd-10;
        fc1_weights[48][186] = 16'sd50;
        fc1_weights[48][187] = 16'sd35;
        fc1_weights[48][188] = 16'sd-14;
        fc1_weights[48][189] = 16'sd21;
        fc1_weights[48][190] = 16'sd-4;
        fc1_weights[48][191] = 16'sd-36;
        fc1_weights[48][192] = 16'sd-18;
        fc1_weights[48][193] = 16'sd-3;
        fc1_weights[48][194] = 16'sd-20;
        fc1_weights[48][195] = 16'sd14;
        fc1_weights[48][196] = 16'sd23;
        fc1_weights[48][197] = 16'sd6;
        fc1_weights[48][198] = 16'sd-12;
        fc1_weights[48][199] = 16'sd18;
        fc1_weights[48][200] = 16'sd7;
        fc1_weights[48][201] = 16'sd8;
        fc1_weights[48][202] = 16'sd-6;
        fc1_weights[48][203] = 16'sd23;
        fc1_weights[48][204] = 16'sd45;
        fc1_weights[48][205] = 16'sd0;
        fc1_weights[48][206] = 16'sd3;
        fc1_weights[48][207] = 16'sd32;
        fc1_weights[49][0] = 16'sd-18;
        fc1_weights[49][1] = 16'sd8;
        fc1_weights[49][2] = 16'sd-24;
        fc1_weights[49][3] = 16'sd-51;
        fc1_weights[49][4] = 16'sd-32;
        fc1_weights[49][5] = 16'sd-27;
        fc1_weights[49][6] = 16'sd-69;
        fc1_weights[49][7] = 16'sd16;
        fc1_weights[49][8] = 16'sd-14;
        fc1_weights[49][9] = 16'sd-34;
        fc1_weights[49][10] = 16'sd17;
        fc1_weights[49][11] = 16'sd64;
        fc1_weights[49][12] = 16'sd-5;
        fc1_weights[49][13] = 16'sd-9;
        fc1_weights[49][14] = 16'sd-26;
        fc1_weights[49][15] = 16'sd-23;
        fc1_weights[49][16] = 16'sd-6;
        fc1_weights[49][17] = 16'sd-7;
        fc1_weights[49][18] = 16'sd2;
        fc1_weights[49][19] = 16'sd-47;
        fc1_weights[49][20] = 16'sd0;
        fc1_weights[49][21] = 16'sd10;
        fc1_weights[49][22] = 16'sd3;
        fc1_weights[49][23] = 16'sd-1;
        fc1_weights[49][24] = 16'sd51;
        fc1_weights[49][25] = 16'sd50;
        fc1_weights[49][26] = 16'sd-7;
        fc1_weights[49][27] = 16'sd-17;
        fc1_weights[49][28] = 16'sd-40;
        fc1_weights[49][29] = 16'sd5;
        fc1_weights[49][30] = 16'sd-8;
        fc1_weights[49][31] = 16'sd-17;
        fc1_weights[49][32] = 16'sd-33;
        fc1_weights[49][33] = 16'sd-51;
        fc1_weights[49][34] = 16'sd32;
        fc1_weights[49][35] = 16'sd25;
        fc1_weights[49][36] = 16'sd54;
        fc1_weights[49][37] = 16'sd12;
        fc1_weights[49][38] = 16'sd8;
        fc1_weights[49][39] = 16'sd-23;
        fc1_weights[49][40] = 16'sd-17;
        fc1_weights[49][41] = 16'sd-4;
        fc1_weights[49][42] = 16'sd-28;
        fc1_weights[49][43] = 16'sd-23;
        fc1_weights[49][44] = 16'sd-11;
        fc1_weights[49][45] = 16'sd-9;
        fc1_weights[49][46] = 16'sd10;
        fc1_weights[49][47] = 16'sd9;
        fc1_weights[49][48] = 16'sd-13;
        fc1_weights[49][49] = 16'sd24;
        fc1_weights[49][50] = 16'sd5;
        fc1_weights[49][51] = 16'sd-1;
        fc1_weights[49][52] = 16'sd-15;
        fc1_weights[49][53] = 16'sd-4;
        fc1_weights[49][54] = 16'sd-9;
        fc1_weights[49][55] = 16'sd5;
        fc1_weights[49][56] = 16'sd21;
        fc1_weights[49][57] = 16'sd38;
        fc1_weights[49][58] = 16'sd-8;
        fc1_weights[49][59] = 16'sd-31;
        fc1_weights[49][60] = 16'sd55;
        fc1_weights[49][61] = 16'sd37;
        fc1_weights[49][62] = 16'sd18;
        fc1_weights[49][63] = 16'sd58;
        fc1_weights[49][64] = 16'sd83;
        fc1_weights[49][65] = 16'sd-28;
        fc1_weights[49][66] = 16'sd2;
        fc1_weights[49][67] = 16'sd12;
        fc1_weights[49][68] = 16'sd-45;
        fc1_weights[49][69] = 16'sd-7;
        fc1_weights[49][70] = 16'sd-1;
        fc1_weights[49][71] = 16'sd-21;
        fc1_weights[49][72] = 16'sd-2;
        fc1_weights[49][73] = 16'sd14;
        fc1_weights[49][74] = 16'sd33;
        fc1_weights[49][75] = 16'sd-8;
        fc1_weights[49][76] = 16'sd-9;
        fc1_weights[49][77] = 16'sd48;
        fc1_weights[49][78] = 16'sd-22;
        fc1_weights[49][79] = 16'sd-51;
        fc1_weights[49][80] = 16'sd-19;
        fc1_weights[49][81] = 16'sd-12;
        fc1_weights[49][82] = 16'sd-3;
        fc1_weights[49][83] = 16'sd-14;
        fc1_weights[49][84] = 16'sd2;
        fc1_weights[49][85] = 16'sd-32;
        fc1_weights[49][86] = 16'sd-27;
        fc1_weights[49][87] = 16'sd35;
        fc1_weights[49][88] = 16'sd37;
        fc1_weights[49][89] = 16'sd-37;
        fc1_weights[49][90] = 16'sd23;
        fc1_weights[49][91] = 16'sd8;
        fc1_weights[49][92] = 16'sd16;
        fc1_weights[49][93] = 16'sd-21;
        fc1_weights[49][94] = 16'sd-19;
        fc1_weights[49][95] = 16'sd-12;
        fc1_weights[49][96] = 16'sd-10;
        fc1_weights[49][97] = 16'sd31;
        fc1_weights[49][98] = 16'sd41;
        fc1_weights[49][99] = 16'sd-1;
        fc1_weights[49][100] = 16'sd31;
        fc1_weights[49][101] = 16'sd28;
        fc1_weights[49][102] = 16'sd4;
        fc1_weights[49][103] = 16'sd26;
        fc1_weights[49][104] = 16'sd7;
        fc1_weights[49][105] = 16'sd-32;
        fc1_weights[49][106] = 16'sd-12;
        fc1_weights[49][107] = 16'sd-14;
        fc1_weights[49][108] = 16'sd14;
        fc1_weights[49][109] = 16'sd-20;
        fc1_weights[49][110] = 16'sd8;
        fc1_weights[49][111] = 16'sd-23;
        fc1_weights[49][112] = 16'sd37;
        fc1_weights[49][113] = 16'sd34;
        fc1_weights[49][114] = 16'sd28;
        fc1_weights[49][115] = 16'sd31;
        fc1_weights[49][116] = 16'sd36;
        fc1_weights[49][117] = 16'sd33;
        fc1_weights[49][118] = 16'sd-11;
        fc1_weights[49][119] = 16'sd-49;
        fc1_weights[49][120] = 16'sd-32;
        fc1_weights[49][121] = 16'sd-13;
        fc1_weights[49][122] = 16'sd-12;
        fc1_weights[49][123] = 16'sd-3;
        fc1_weights[49][124] = 16'sd-20;
        fc1_weights[49][125] = 16'sd21;
        fc1_weights[49][126] = 16'sd43;
        fc1_weights[49][127] = 16'sd14;
        fc1_weights[49][128] = 16'sd1;
        fc1_weights[49][129] = 16'sd15;
        fc1_weights[49][130] = 16'sd-41;
        fc1_weights[49][131] = 16'sd-4;
        fc1_weights[49][132] = 16'sd9;
        fc1_weights[49][133] = 16'sd-15;
        fc1_weights[49][134] = 16'sd-4;
        fc1_weights[49][135] = 16'sd-29;
        fc1_weights[49][136] = 16'sd-2;
        fc1_weights[49][137] = 16'sd-47;
        fc1_weights[49][138] = 16'sd71;
        fc1_weights[49][139] = 16'sd2;
        fc1_weights[49][140] = 16'sd-3;
        fc1_weights[49][141] = 16'sd20;
        fc1_weights[49][142] = 16'sd-20;
        fc1_weights[49][143] = 16'sd23;
        fc1_weights[49][144] = 16'sd34;
        fc1_weights[49][145] = 16'sd18;
        fc1_weights[49][146] = 16'sd15;
        fc1_weights[49][147] = 16'sd0;
        fc1_weights[49][148] = 16'sd-5;
        fc1_weights[49][149] = 16'sd34;
        fc1_weights[49][150] = 16'sd26;
        fc1_weights[49][151] = 16'sd76;
        fc1_weights[49][152] = 16'sd-15;
        fc1_weights[49][153] = 16'sd18;
        fc1_weights[49][154] = 16'sd18;
        fc1_weights[49][155] = 16'sd33;
        fc1_weights[49][156] = 16'sd-20;
        fc1_weights[49][157] = 16'sd-24;
        fc1_weights[49][158] = 16'sd-25;
        fc1_weights[49][159] = 16'sd20;
        fc1_weights[49][160] = 16'sd-15;
        fc1_weights[49][161] = 16'sd6;
        fc1_weights[49][162] = 16'sd45;
        fc1_weights[49][163] = 16'sd-41;
        fc1_weights[49][164] = 16'sd-27;
        fc1_weights[49][165] = 16'sd-20;
        fc1_weights[49][166] = 16'sd-29;
        fc1_weights[49][167] = 16'sd17;
        fc1_weights[49][168] = 16'sd15;
        fc1_weights[49][169] = 16'sd9;
        fc1_weights[49][170] = 16'sd49;
        fc1_weights[49][171] = 16'sd-42;
        fc1_weights[49][172] = 16'sd14;
        fc1_weights[49][173] = 16'sd16;
        fc1_weights[49][174] = 16'sd-1;
        fc1_weights[49][175] = 16'sd2;
        fc1_weights[49][176] = 16'sd-7;
        fc1_weights[49][177] = 16'sd9;
        fc1_weights[49][178] = 16'sd20;
        fc1_weights[49][179] = 16'sd40;
        fc1_weights[49][180] = 16'sd1;
        fc1_weights[49][181] = 16'sd10;
        fc1_weights[49][182] = 16'sd7;
        fc1_weights[49][183] = 16'sd-19;
        fc1_weights[49][184] = 16'sd-7;
        fc1_weights[49][185] = 16'sd19;
        fc1_weights[49][186] = 16'sd11;
        fc1_weights[49][187] = 16'sd-29;
        fc1_weights[49][188] = 16'sd-8;
        fc1_weights[49][189] = 16'sd-53;
        fc1_weights[49][190] = 16'sd13;
        fc1_weights[49][191] = 16'sd-4;
        fc1_weights[49][192] = 16'sd-5;
        fc1_weights[49][193] = 16'sd-13;
        fc1_weights[49][194] = 16'sd-33;
        fc1_weights[49][195] = 16'sd13;
        fc1_weights[49][196] = 16'sd1;
        fc1_weights[49][197] = 16'sd15;
        fc1_weights[49][198] = 16'sd-40;
        fc1_weights[49][199] = 16'sd-24;
        fc1_weights[49][200] = 16'sd18;
        fc1_weights[49][201] = 16'sd-44;
        fc1_weights[49][202] = 16'sd-64;
        fc1_weights[49][203] = 16'sd39;
        fc1_weights[49][204] = 16'sd-13;
        fc1_weights[49][205] = 16'sd8;
        fc1_weights[49][206] = 16'sd-17;
        fc1_weights[49][207] = 16'sd36;
        fc1_weights[50][0] = 16'sd44;
        fc1_weights[50][1] = 16'sd23;
        fc1_weights[50][2] = 16'sd2;
        fc1_weights[50][3] = 16'sd14;
        fc1_weights[50][4] = 16'sd35;
        fc1_weights[50][5] = 16'sd30;
        fc1_weights[50][6] = 16'sd8;
        fc1_weights[50][7] = 16'sd14;
        fc1_weights[50][8] = 16'sd5;
        fc1_weights[50][9] = 16'sd20;
        fc1_weights[50][10] = 16'sd-48;
        fc1_weights[50][11] = 16'sd-6;
        fc1_weights[50][12] = 16'sd2;
        fc1_weights[50][13] = 16'sd-6;
        fc1_weights[50][14] = 16'sd3;
        fc1_weights[50][15] = 16'sd10;
        fc1_weights[50][16] = 16'sd-17;
        fc1_weights[50][17] = 16'sd-1;
        fc1_weights[50][18] = 16'sd3;
        fc1_weights[50][19] = 16'sd5;
        fc1_weights[50][20] = 16'sd16;
        fc1_weights[50][21] = 16'sd2;
        fc1_weights[50][22] = 16'sd1;
        fc1_weights[50][23] = 16'sd39;
        fc1_weights[50][24] = 16'sd37;
        fc1_weights[50][25] = 16'sd-2;
        fc1_weights[50][26] = 16'sd4;
        fc1_weights[50][27] = 16'sd25;
        fc1_weights[50][28] = 16'sd17;
        fc1_weights[50][29] = 16'sd14;
        fc1_weights[50][30] = 16'sd23;
        fc1_weights[50][31] = 16'sd48;
        fc1_weights[50][32] = 16'sd35;
        fc1_weights[50][33] = 16'sd26;
        fc1_weights[50][34] = 16'sd-35;
        fc1_weights[50][35] = 16'sd11;
        fc1_weights[50][36] = 16'sd-4;
        fc1_weights[50][37] = 16'sd8;
        fc1_weights[50][38] = 16'sd18;
        fc1_weights[50][39] = 16'sd12;
        fc1_weights[50][40] = 16'sd-16;
        fc1_weights[50][41] = 16'sd-10;
        fc1_weights[50][42] = 16'sd14;
        fc1_weights[50][43] = 16'sd-20;
        fc1_weights[50][44] = 16'sd-13;
        fc1_weights[50][45] = 16'sd-27;
        fc1_weights[50][46] = 16'sd-6;
        fc1_weights[50][47] = 16'sd-15;
        fc1_weights[50][48] = 16'sd-10;
        fc1_weights[50][49] = 16'sd-22;
        fc1_weights[50][50] = 16'sd-28;
        fc1_weights[50][51] = 16'sd-12;
        fc1_weights[50][52] = 16'sd-3;
        fc1_weights[50][53] = 16'sd19;
        fc1_weights[50][54] = 16'sd24;
        fc1_weights[50][55] = 16'sd16;
        fc1_weights[50][56] = 16'sd28;
        fc1_weights[50][57] = 16'sd33;
        fc1_weights[50][58] = 16'sd27;
        fc1_weights[50][59] = 16'sd16;
        fc1_weights[50][60] = 16'sd7;
        fc1_weights[50][61] = 16'sd29;
        fc1_weights[50][62] = 16'sd0;
        fc1_weights[50][63] = 16'sd5;
        fc1_weights[50][64] = 16'sd35;
        fc1_weights[50][65] = 16'sd-33;
        fc1_weights[50][66] = 16'sd-41;
        fc1_weights[50][67] = 16'sd-34;
        fc1_weights[50][68] = 16'sd-22;
        fc1_weights[50][69] = 16'sd-10;
        fc1_weights[50][70] = 16'sd-32;
        fc1_weights[50][71] = 16'sd22;
        fc1_weights[50][72] = 16'sd36;
        fc1_weights[50][73] = 16'sd-15;
        fc1_weights[50][74] = 16'sd-5;
        fc1_weights[50][75] = 16'sd-31;
        fc1_weights[50][76] = 16'sd-27;
        fc1_weights[50][77] = 16'sd-6;
        fc1_weights[50][78] = 16'sd30;
        fc1_weights[50][79] = 16'sd32;
        fc1_weights[50][80] = 16'sd29;
        fc1_weights[50][81] = 16'sd-4;
        fc1_weights[50][82] = 16'sd32;
        fc1_weights[50][83] = 16'sd5;
        fc1_weights[50][84] = 16'sd24;
        fc1_weights[50][85] = 16'sd39;
        fc1_weights[50][86] = 16'sd30;
        fc1_weights[50][87] = 16'sd22;
        fc1_weights[50][88] = 16'sd-13;
        fc1_weights[50][89] = 16'sd-3;
        fc1_weights[50][90] = 16'sd33;
        fc1_weights[50][91] = 16'sd0;
        fc1_weights[50][92] = 16'sd-24;
        fc1_weights[50][93] = 16'sd-17;
        fc1_weights[50][94] = 16'sd-13;
        fc1_weights[50][95] = 16'sd8;
        fc1_weights[50][96] = 16'sd-41;
        fc1_weights[50][97] = 16'sd-27;
        fc1_weights[50][98] = 16'sd3;
        fc1_weights[50][99] = 16'sd-20;
        fc1_weights[50][100] = 16'sd18;
        fc1_weights[50][101] = 16'sd-27;
        fc1_weights[50][102] = 16'sd-30;
        fc1_weights[50][103] = 16'sd-14;
        fc1_weights[50][104] = 16'sd3;
        fc1_weights[50][105] = 16'sd11;
        fc1_weights[50][106] = 16'sd32;
        fc1_weights[50][107] = 16'sd4;
        fc1_weights[50][108] = 16'sd-1;
        fc1_weights[50][109] = 16'sd-9;
        fc1_weights[50][110] = 16'sd-1;
        fc1_weights[50][111] = 16'sd-28;
        fc1_weights[50][112] = 16'sd4;
        fc1_weights[50][113] = 16'sd26;
        fc1_weights[50][114] = 16'sd6;
        fc1_weights[50][115] = 16'sd-35;
        fc1_weights[50][116] = 16'sd50;
        fc1_weights[50][117] = 16'sd-9;
        fc1_weights[50][118] = 16'sd-5;
        fc1_weights[50][119] = 16'sd3;
        fc1_weights[50][120] = 16'sd-6;
        fc1_weights[50][121] = 16'sd-13;
        fc1_weights[50][122] = 16'sd-45;
        fc1_weights[50][123] = 16'sd11;
        fc1_weights[50][124] = 16'sd-9;
        fc1_weights[50][125] = 16'sd27;
        fc1_weights[50][126] = 16'sd-18;
        fc1_weights[50][127] = 16'sd-34;
        fc1_weights[50][128] = 16'sd-23;
        fc1_weights[50][129] = 16'sd-33;
        fc1_weights[50][130] = 16'sd-15;
        fc1_weights[50][131] = 16'sd-18;
        fc1_weights[50][132] = 16'sd-9;
        fc1_weights[50][133] = 16'sd-18;
        fc1_weights[50][134] = 16'sd-12;
        fc1_weights[50][135] = 16'sd-42;
        fc1_weights[50][136] = 16'sd-42;
        fc1_weights[50][137] = 16'sd18;
        fc1_weights[50][138] = 16'sd19;
        fc1_weights[50][139] = 16'sd-6;
        fc1_weights[50][140] = 16'sd2;
        fc1_weights[50][141] = 16'sd-53;
        fc1_weights[50][142] = 16'sd-5;
        fc1_weights[50][143] = 16'sd24;
        fc1_weights[50][144] = 16'sd-23;
        fc1_weights[50][145] = 16'sd-33;
        fc1_weights[50][146] = 16'sd-28;
        fc1_weights[50][147] = 16'sd-11;
        fc1_weights[50][148] = 16'sd-21;
        fc1_weights[50][149] = 16'sd-39;
        fc1_weights[50][150] = 16'sd-46;
        fc1_weights[50][151] = 16'sd7;
        fc1_weights[50][152] = 16'sd-13;
        fc1_weights[50][153] = 16'sd9;
        fc1_weights[50][154] = 16'sd-7;
        fc1_weights[50][155] = 16'sd53;
        fc1_weights[50][156] = 16'sd7;
        fc1_weights[50][157] = 16'sd-2;
        fc1_weights[50][158] = 16'sd-15;
        fc1_weights[50][159] = 16'sd-37;
        fc1_weights[50][160] = 16'sd-47;
        fc1_weights[50][161] = 16'sd-25;
        fc1_weights[50][162] = 16'sd0;
        fc1_weights[50][163] = 16'sd5;
        fc1_weights[50][164] = 16'sd10;
        fc1_weights[50][165] = 16'sd-29;
        fc1_weights[50][166] = 16'sd23;
        fc1_weights[50][167] = 16'sd9;
        fc1_weights[50][168] = 16'sd3;
        fc1_weights[50][169] = 16'sd15;
        fc1_weights[50][170] = 16'sd4;
        fc1_weights[50][171] = 16'sd2;
        fc1_weights[50][172] = 16'sd-25;
        fc1_weights[50][173] = 16'sd-13;
        fc1_weights[50][174] = 16'sd12;
        fc1_weights[50][175] = 16'sd25;
        fc1_weights[50][176] = 16'sd22;
        fc1_weights[50][177] = 16'sd-17;
        fc1_weights[50][178] = 16'sd-39;
        fc1_weights[50][179] = 16'sd24;
        fc1_weights[50][180] = 16'sd-21;
        fc1_weights[50][181] = 16'sd3;
        fc1_weights[50][182] = 16'sd-34;
        fc1_weights[50][183] = 16'sd-25;
        fc1_weights[50][184] = 16'sd-25;
        fc1_weights[50][185] = 16'sd-12;
        fc1_weights[50][186] = 16'sd-27;
        fc1_weights[50][187] = 16'sd-7;
        fc1_weights[50][188] = 16'sd-34;
        fc1_weights[50][189] = 16'sd-6;
        fc1_weights[50][190] = 16'sd15;
        fc1_weights[50][191] = 16'sd6;
        fc1_weights[50][192] = 16'sd-2;
        fc1_weights[50][193] = 16'sd12;
        fc1_weights[50][194] = 16'sd31;
        fc1_weights[50][195] = 16'sd-14;
        fc1_weights[50][196] = 16'sd19;
        fc1_weights[50][197] = 16'sd-9;
        fc1_weights[50][198] = 16'sd-2;
        fc1_weights[50][199] = 16'sd17;
        fc1_weights[50][200] = 16'sd4;
        fc1_weights[50][201] = 16'sd0;
        fc1_weights[50][202] = 16'sd-2;
        fc1_weights[50][203] = 16'sd7;
        fc1_weights[50][204] = 16'sd-7;
        fc1_weights[50][205] = 16'sd-9;
        fc1_weights[50][206] = 16'sd-19;
        fc1_weights[50][207] = 16'sd-27;
        fc1_weights[51][0] = 16'sd-25;
        fc1_weights[51][1] = 16'sd23;
        fc1_weights[51][2] = 16'sd8;
        fc1_weights[51][3] = 16'sd-31;
        fc1_weights[51][4] = 16'sd4;
        fc1_weights[51][5] = 16'sd38;
        fc1_weights[51][6] = 16'sd37;
        fc1_weights[51][7] = 16'sd62;
        fc1_weights[51][8] = 16'sd59;
        fc1_weights[51][9] = 16'sd51;
        fc1_weights[51][10] = 16'sd-1;
        fc1_weights[51][11] = 16'sd30;
        fc1_weights[51][12] = 16'sd11;
        fc1_weights[51][13] = 16'sd-23;
        fc1_weights[51][14] = 16'sd-76;
        fc1_weights[51][15] = 16'sd-14;
        fc1_weights[51][16] = 16'sd-35;
        fc1_weights[51][17] = 16'sd-28;
        fc1_weights[51][18] = 16'sd-2;
        fc1_weights[51][19] = 16'sd-61;
        fc1_weights[51][20] = 16'sd8;
        fc1_weights[51][21] = 16'sd-39;
        fc1_weights[51][22] = 16'sd0;
        fc1_weights[51][23] = 16'sd47;
        fc1_weights[51][24] = 16'sd23;
        fc1_weights[51][25] = 16'sd12;
        fc1_weights[51][26] = 16'sd-6;
        fc1_weights[51][27] = 16'sd-17;
        fc1_weights[51][28] = 16'sd-11;
        fc1_weights[51][29] = 16'sd14;
        fc1_weights[51][30] = 16'sd32;
        fc1_weights[51][31] = 16'sd87;
        fc1_weights[51][32] = 16'sd3;
        fc1_weights[51][33] = 16'sd-52;
        fc1_weights[51][34] = 16'sd61;
        fc1_weights[51][35] = 16'sd44;
        fc1_weights[51][36] = 16'sd85;
        fc1_weights[51][37] = 16'sd-44;
        fc1_weights[51][38] = 16'sd0;
        fc1_weights[51][39] = 16'sd12;
        fc1_weights[51][40] = 16'sd-28;
        fc1_weights[51][41] = 16'sd-81;
        fc1_weights[51][42] = 16'sd-24;
        fc1_weights[51][43] = 16'sd-61;
        fc1_weights[51][44] = 16'sd-17;
        fc1_weights[51][45] = 16'sd26;
        fc1_weights[51][46] = 16'sd-45;
        fc1_weights[51][47] = 16'sd2;
        fc1_weights[51][48] = 16'sd10;
        fc1_weights[51][49] = 16'sd66;
        fc1_weights[51][50] = 16'sd-40;
        fc1_weights[51][51] = 16'sd11;
        fc1_weights[51][52] = 16'sd45;
        fc1_weights[51][53] = 16'sd-30;
        fc1_weights[51][54] = 16'sd-38;
        fc1_weights[51][55] = 16'sd-79;
        fc1_weights[51][56] = 16'sd9;
        fc1_weights[51][57] = 16'sd-24;
        fc1_weights[51][58] = 16'sd-32;
        fc1_weights[51][59] = 16'sd9;
        fc1_weights[51][60] = 16'sd84;
        fc1_weights[51][61] = 16'sd-16;
        fc1_weights[51][62] = 16'sd-20;
        fc1_weights[51][63] = 16'sd1;
        fc1_weights[51][64] = 16'sd93;
        fc1_weights[51][65] = 16'sd-19;
        fc1_weights[51][66] = 16'sd82;
        fc1_weights[51][67] = 16'sd-9;
        fc1_weights[51][68] = 16'sd-76;
        fc1_weights[51][69] = 16'sd17;
        fc1_weights[51][70] = 16'sd56;
        fc1_weights[51][71] = 16'sd122;
        fc1_weights[51][72] = 16'sd49;
        fc1_weights[51][73] = 16'sd25;
        fc1_weights[51][74] = 16'sd67;
        fc1_weights[51][75] = 16'sd-5;
        fc1_weights[51][76] = 16'sd41;
        fc1_weights[51][77] = 16'sd35;
        fc1_weights[51][78] = 16'sd74;
        fc1_weights[51][79] = 16'sd106;
        fc1_weights[51][80] = 16'sd-29;
        fc1_weights[51][81] = 16'sd6;
        fc1_weights[51][82] = 16'sd11;
        fc1_weights[51][83] = 16'sd68;
        fc1_weights[51][84] = 16'sd-64;
        fc1_weights[51][85] = 16'sd-33;
        fc1_weights[51][86] = 16'sd36;
        fc1_weights[51][87] = 16'sd95;
        fc1_weights[51][88] = 16'sd43;
        fc1_weights[51][89] = 16'sd-12;
        fc1_weights[51][90] = 16'sd49;
        fc1_weights[51][91] = 16'sd34;
        fc1_weights[51][92] = 16'sd-14;
        fc1_weights[51][93] = 16'sd-64;
        fc1_weights[51][94] = 16'sd-109;
        fc1_weights[51][95] = 16'sd42;
        fc1_weights[51][96] = 16'sd-18;
        fc1_weights[51][97] = 16'sd21;
        fc1_weights[51][98] = 16'sd-41;
        fc1_weights[51][99] = 16'sd-65;
        fc1_weights[51][100] = 16'sd-18;
        fc1_weights[51][101] = 16'sd-53;
        fc1_weights[51][102] = 16'sd-56;
        fc1_weights[51][103] = 16'sd25;
        fc1_weights[51][104] = 16'sd97;
        fc1_weights[51][105] = 16'sd4;
        fc1_weights[51][106] = 16'sd48;
        fc1_weights[51][107] = 16'sd77;
        fc1_weights[51][108] = 16'sd-19;
        fc1_weights[51][109] = 16'sd44;
        fc1_weights[51][110] = 16'sd-39;
        fc1_weights[51][111] = 16'sd28;
        fc1_weights[51][112] = 16'sd101;
        fc1_weights[51][113] = 16'sd-14;
        fc1_weights[51][114] = 16'sd9;
        fc1_weights[51][115] = 16'sd-9;
        fc1_weights[51][116] = 16'sd8;
        fc1_weights[51][117] = 16'sd43;
        fc1_weights[51][118] = 16'sd21;
        fc1_weights[51][119] = 16'sd2;
        fc1_weights[51][120] = 16'sd-30;
        fc1_weights[51][121] = 16'sd78;
        fc1_weights[51][122] = 16'sd25;
        fc1_weights[51][123] = 16'sd122;
        fc1_weights[51][124] = 16'sd8;
        fc1_weights[51][125] = 16'sd-24;
        fc1_weights[51][126] = 16'sd-11;
        fc1_weights[51][127] = 16'sd-9;
        fc1_weights[51][128] = 16'sd23;
        fc1_weights[51][129] = 16'sd34;
        fc1_weights[51][130] = 16'sd49;
        fc1_weights[51][131] = 16'sd82;
        fc1_weights[51][132] = 16'sd9;
        fc1_weights[51][133] = 16'sd46;
        fc1_weights[51][134] = 16'sd-19;
        fc1_weights[51][135] = 16'sd11;
        fc1_weights[51][136] = 16'sd-30;
        fc1_weights[51][137] = 16'sd-6;
        fc1_weights[51][138] = 16'sd-14;
        fc1_weights[51][139] = 16'sd-111;
        fc1_weights[51][140] = 16'sd-72;
        fc1_weights[51][141] = 16'sd-35;
        fc1_weights[51][142] = 16'sd72;
        fc1_weights[51][143] = 16'sd-14;
        fc1_weights[51][144] = 16'sd62;
        fc1_weights[51][145] = 16'sd-5;
        fc1_weights[51][146] = 16'sd14;
        fc1_weights[51][147] = 16'sd-43;
        fc1_weights[51][148] = 16'sd20;
        fc1_weights[51][149] = 16'sd-21;
        fc1_weights[51][150] = 16'sd-3;
        fc1_weights[51][151] = 16'sd-21;
        fc1_weights[51][152] = 16'sd-32;
        fc1_weights[51][153] = 16'sd-48;
        fc1_weights[51][154] = 16'sd2;
        fc1_weights[51][155] = 16'sd20;
        fc1_weights[51][156] = 16'sd44;
        fc1_weights[51][157] = 16'sd20;
        fc1_weights[51][158] = 16'sd-63;
        fc1_weights[51][159] = 16'sd-26;
        fc1_weights[51][160] = 16'sd-16;
        fc1_weights[51][161] = 16'sd8;
        fc1_weights[51][162] = 16'sd3;
        fc1_weights[51][163] = 16'sd-6;
        fc1_weights[51][164] = 16'sd-62;
        fc1_weights[51][165] = 16'sd-52;
        fc1_weights[51][166] = 16'sd-21;
        fc1_weights[51][167] = 16'sd-28;
        fc1_weights[51][168] = 16'sd-22;
        fc1_weights[51][169] = 16'sd11;
        fc1_weights[51][170] = 16'sd24;
        fc1_weights[51][171] = 16'sd2;
        fc1_weights[51][172] = 16'sd-37;
        fc1_weights[51][173] = 16'sd-5;
        fc1_weights[51][174] = 16'sd25;
        fc1_weights[51][175] = 16'sd-21;
        fc1_weights[51][176] = 16'sd-39;
        fc1_weights[51][177] = 16'sd20;
        fc1_weights[51][178] = 16'sd-8;
        fc1_weights[51][179] = 16'sd-4;
        fc1_weights[51][180] = 16'sd20;
        fc1_weights[51][181] = 16'sd11;
        fc1_weights[51][182] = 16'sd16;
        fc1_weights[51][183] = 16'sd21;
        fc1_weights[51][184] = 16'sd-1;
        fc1_weights[51][185] = 16'sd-11;
        fc1_weights[51][186] = 16'sd-32;
        fc1_weights[51][187] = 16'sd-40;
        fc1_weights[51][188] = 16'sd-18;
        fc1_weights[51][189] = 16'sd-16;
        fc1_weights[51][190] = 16'sd-56;
        fc1_weights[51][191] = 16'sd14;
        fc1_weights[51][192] = 16'sd-14;
        fc1_weights[51][193] = 16'sd-39;
        fc1_weights[51][194] = 16'sd7;
        fc1_weights[51][195] = 16'sd-17;
        fc1_weights[51][196] = 16'sd6;
        fc1_weights[51][197] = 16'sd42;
        fc1_weights[51][198] = 16'sd-14;
        fc1_weights[51][199] = 16'sd-43;
        fc1_weights[51][200] = 16'sd12;
        fc1_weights[51][201] = 16'sd-1;
        fc1_weights[51][202] = 16'sd-13;
        fc1_weights[51][203] = 16'sd-11;
        fc1_weights[51][204] = 16'sd-26;
        fc1_weights[51][205] = 16'sd-54;
        fc1_weights[51][206] = 16'sd39;
        fc1_weights[51][207] = 16'sd-10;
        fc1_weights[52][0] = 16'sd41;
        fc1_weights[52][1] = 16'sd-21;
        fc1_weights[52][2] = 16'sd9;
        fc1_weights[52][3] = 16'sd41;
        fc1_weights[52][4] = 16'sd27;
        fc1_weights[52][5] = 16'sd67;
        fc1_weights[52][6] = 16'sd12;
        fc1_weights[52][7] = 16'sd31;
        fc1_weights[52][8] = 16'sd6;
        fc1_weights[52][9] = 16'sd28;
        fc1_weights[52][10] = 16'sd-4;
        fc1_weights[52][11] = 16'sd92;
        fc1_weights[52][12] = 16'sd-45;
        fc1_weights[52][13] = 16'sd37;
        fc1_weights[52][14] = 16'sd-1;
        fc1_weights[52][15] = 16'sd3;
        fc1_weights[52][16] = 16'sd-43;
        fc1_weights[52][17] = 16'sd-30;
        fc1_weights[52][18] = 16'sd38;
        fc1_weights[52][19] = 16'sd-21;
        fc1_weights[52][20] = 16'sd-8;
        fc1_weights[52][21] = 16'sd-21;
        fc1_weights[52][22] = 16'sd16;
        fc1_weights[52][23] = 16'sd-31;
        fc1_weights[52][24] = 16'sd7;
        fc1_weights[52][25] = 16'sd-28;
        fc1_weights[52][26] = 16'sd-35;
        fc1_weights[52][27] = 16'sd-9;
        fc1_weights[52][28] = 16'sd-61;
        fc1_weights[52][29] = 16'sd-5;
        fc1_weights[52][30] = 16'sd13;
        fc1_weights[52][31] = 16'sd80;
        fc1_weights[52][32] = 16'sd31;
        fc1_weights[52][33] = 16'sd54;
        fc1_weights[52][34] = 16'sd39;
        fc1_weights[52][35] = 16'sd13;
        fc1_weights[52][36] = 16'sd17;
        fc1_weights[52][37] = 16'sd22;
        fc1_weights[52][38] = 16'sd-13;
        fc1_weights[52][39] = 16'sd-112;
        fc1_weights[52][40] = 16'sd26;
        fc1_weights[52][41] = 16'sd-31;
        fc1_weights[52][42] = 16'sd9;
        fc1_weights[52][43] = 16'sd76;
        fc1_weights[52][44] = 16'sd19;
        fc1_weights[52][45] = 16'sd-20;
        fc1_weights[52][46] = 16'sd36;
        fc1_weights[52][47] = 16'sd21;
        fc1_weights[52][48] = 16'sd-16;
        fc1_weights[52][49] = 16'sd-3;
        fc1_weights[52][50] = 16'sd-42;
        fc1_weights[52][51] = 16'sd-30;
        fc1_weights[52][52] = 16'sd-35;
        fc1_weights[52][53] = 16'sd42;
        fc1_weights[52][54] = 16'sd-59;
        fc1_weights[52][55] = 16'sd6;
        fc1_weights[52][56] = 16'sd0;
        fc1_weights[52][57] = 16'sd79;
        fc1_weights[52][58] = 16'sd80;
        fc1_weights[52][59] = 16'sd29;
        fc1_weights[52][60] = 16'sd53;
        fc1_weights[52][61] = 16'sd47;
        fc1_weights[52][62] = 16'sd32;
        fc1_weights[52][63] = 16'sd64;
        fc1_weights[52][64] = 16'sd-70;
        fc1_weights[52][65] = 16'sd-18;
        fc1_weights[52][66] = 16'sd-25;
        fc1_weights[52][67] = 16'sd0;
        fc1_weights[52][68] = 16'sd41;
        fc1_weights[52][69] = 16'sd12;
        fc1_weights[52][70] = 16'sd6;
        fc1_weights[52][71] = 16'sd-41;
        fc1_weights[52][72] = 16'sd23;
        fc1_weights[52][73] = 16'sd29;
        fc1_weights[52][74] = 16'sd-44;
        fc1_weights[52][75] = 16'sd-12;
        fc1_weights[52][76] = 16'sd44;
        fc1_weights[52][77] = 16'sd-10;
        fc1_weights[52][78] = 16'sd-10;
        fc1_weights[52][79] = 16'sd32;
        fc1_weights[52][80] = 16'sd-26;
        fc1_weights[52][81] = 16'sd-41;
        fc1_weights[52][82] = 16'sd-4;
        fc1_weights[52][83] = 16'sd-19;
        fc1_weights[52][84] = 16'sd-5;
        fc1_weights[52][85] = 16'sd-4;
        fc1_weights[52][86] = 16'sd-20;
        fc1_weights[52][87] = 16'sd-16;
        fc1_weights[52][88] = 16'sd-75;
        fc1_weights[52][89] = 16'sd28;
        fc1_weights[52][90] = 16'sd-11;
        fc1_weights[52][91] = 16'sd-57;
        fc1_weights[52][92] = 16'sd-86;
        fc1_weights[52][93] = 16'sd-42;
        fc1_weights[52][94] = 16'sd-20;
        fc1_weights[52][95] = 16'sd7;
        fc1_weights[52][96] = 16'sd-30;
        fc1_weights[52][97] = 16'sd-67;
        fc1_weights[52][98] = 16'sd-34;
        fc1_weights[52][99] = 16'sd8;
        fc1_weights[52][100] = 16'sd-26;
        fc1_weights[52][101] = 16'sd-6;
        fc1_weights[52][102] = 16'sd-48;
        fc1_weights[52][103] = 16'sd-34;
        fc1_weights[52][104] = 16'sd-17;
        fc1_weights[52][105] = 16'sd-59;
        fc1_weights[52][106] = 16'sd-25;
        fc1_weights[52][107] = 16'sd-17;
        fc1_weights[52][108] = 16'sd35;
        fc1_weights[52][109] = 16'sd35;
        fc1_weights[52][110] = 16'sd47;
        fc1_weights[52][111] = 16'sd-26;
        fc1_weights[52][112] = 16'sd11;
        fc1_weights[52][113] = 16'sd22;
        fc1_weights[52][114] = 16'sd47;
        fc1_weights[52][115] = 16'sd36;
        fc1_weights[52][116] = 16'sd39;
        fc1_weights[52][117] = 16'sd12;
        fc1_weights[52][118] = 16'sd-38;
        fc1_weights[52][119] = 16'sd16;
        fc1_weights[52][120] = 16'sd-14;
        fc1_weights[52][121] = 16'sd-14;
        fc1_weights[52][122] = 16'sd-15;
        fc1_weights[52][123] = 16'sd-78;
        fc1_weights[52][124] = 16'sd-37;
        fc1_weights[52][125] = 16'sd-25;
        fc1_weights[52][126] = 16'sd-69;
        fc1_weights[52][127] = 16'sd-51;
        fc1_weights[52][128] = 16'sd-33;
        fc1_weights[52][129] = 16'sd-72;
        fc1_weights[52][130] = 16'sd69;
        fc1_weights[52][131] = 16'sd43;
        fc1_weights[52][132] = 16'sd8;
        fc1_weights[52][133] = 16'sd19;
        fc1_weights[52][134] = 16'sd-5;
        fc1_weights[52][135] = 16'sd9;
        fc1_weights[52][136] = 16'sd-1;
        fc1_weights[52][137] = 16'sd20;
        fc1_weights[52][138] = 16'sd-23;
        fc1_weights[52][139] = 16'sd1;
        fc1_weights[52][140] = 16'sd6;
        fc1_weights[52][141] = 16'sd-39;
        fc1_weights[52][142] = 16'sd-4;
        fc1_weights[52][143] = 16'sd30;
        fc1_weights[52][144] = 16'sd3;
        fc1_weights[52][145] = 16'sd-41;
        fc1_weights[52][146] = 16'sd-33;
        fc1_weights[52][147] = 16'sd18;
        fc1_weights[52][148] = 16'sd-44;
        fc1_weights[52][149] = 16'sd-4;
        fc1_weights[52][150] = 16'sd-57;
        fc1_weights[52][151] = 16'sd-5;
        fc1_weights[52][152] = 16'sd-6;
        fc1_weights[52][153] = 16'sd-22;
        fc1_weights[52][154] = 16'sd17;
        fc1_weights[52][155] = 16'sd64;
        fc1_weights[52][156] = 16'sd-2;
        fc1_weights[52][157] = 16'sd-24;
        fc1_weights[52][158] = 16'sd-7;
        fc1_weights[52][159] = 16'sd18;
        fc1_weights[52][160] = 16'sd-78;
        fc1_weights[52][161] = 16'sd-24;
        fc1_weights[52][162] = 16'sd-6;
        fc1_weights[52][163] = 16'sd-30;
        fc1_weights[52][164] = 16'sd-6;
        fc1_weights[52][165] = 16'sd25;
        fc1_weights[52][166] = 16'sd22;
        fc1_weights[52][167] = 16'sd-19;
        fc1_weights[52][168] = 16'sd-2;
        fc1_weights[52][169] = 16'sd-22;
        fc1_weights[52][170] = 16'sd-7;
        fc1_weights[52][171] = 16'sd3;
        fc1_weights[52][172] = 16'sd15;
        fc1_weights[52][173] = 16'sd-3;
        fc1_weights[52][174] = 16'sd13;
        fc1_weights[52][175] = 16'sd67;
        fc1_weights[52][176] = 16'sd61;
        fc1_weights[52][177] = 16'sd22;
        fc1_weights[52][178] = 16'sd-13;
        fc1_weights[52][179] = 16'sd73;
        fc1_weights[52][180] = 16'sd23;
        fc1_weights[52][181] = 16'sd-16;
        fc1_weights[52][182] = 16'sd-3;
        fc1_weights[52][183] = 16'sd-52;
        fc1_weights[52][184] = 16'sd-15;
        fc1_weights[52][185] = 16'sd51;
        fc1_weights[52][186] = 16'sd-100;
        fc1_weights[52][187] = 16'sd-82;
        fc1_weights[52][188] = 16'sd-28;
        fc1_weights[52][189] = 16'sd-60;
        fc1_weights[52][190] = 16'sd25;
        fc1_weights[52][191] = 16'sd-31;
        fc1_weights[52][192] = 16'sd-52;
        fc1_weights[52][193] = 16'sd-13;
        fc1_weights[52][194] = 16'sd-43;
        fc1_weights[52][195] = 16'sd-38;
        fc1_weights[52][196] = 16'sd-39;
        fc1_weights[52][197] = 16'sd-5;
        fc1_weights[52][198] = 16'sd-31;
        fc1_weights[52][199] = 16'sd18;
        fc1_weights[52][200] = 16'sd-27;
        fc1_weights[52][201] = 16'sd-9;
        fc1_weights[52][202] = 16'sd0;
        fc1_weights[52][203] = 16'sd71;
        fc1_weights[52][204] = 16'sd16;
        fc1_weights[52][205] = 16'sd54;
        fc1_weights[52][206] = 16'sd-25;
        fc1_weights[52][207] = 16'sd7;
        fc1_weights[53][0] = 16'sd6;
        fc1_weights[53][1] = 16'sd20;
        fc1_weights[53][2] = 16'sd52;
        fc1_weights[53][3] = 16'sd16;
        fc1_weights[53][4] = 16'sd29;
        fc1_weights[53][5] = 16'sd12;
        fc1_weights[53][6] = 16'sd13;
        fc1_weights[53][7] = 16'sd36;
        fc1_weights[53][8] = 16'sd30;
        fc1_weights[53][9] = 16'sd-7;
        fc1_weights[53][10] = 16'sd24;
        fc1_weights[53][11] = 16'sd-10;
        fc1_weights[53][12] = 16'sd-9;
        fc1_weights[53][13] = 16'sd35;
        fc1_weights[53][14] = 16'sd9;
        fc1_weights[53][15] = 16'sd-14;
        fc1_weights[53][16] = 16'sd-10;
        fc1_weights[53][17] = 16'sd61;
        fc1_weights[53][18] = 16'sd35;
        fc1_weights[53][19] = 16'sd1;
        fc1_weights[53][20] = 16'sd-12;
        fc1_weights[53][21] = 16'sd64;
        fc1_weights[53][22] = 16'sd42;
        fc1_weights[53][23] = 16'sd74;
        fc1_weights[53][24] = 16'sd61;
        fc1_weights[53][25] = 16'sd67;
        fc1_weights[53][26] = 16'sd-1;
        fc1_weights[53][27] = 16'sd15;
        fc1_weights[53][28] = 16'sd70;
        fc1_weights[53][29] = 16'sd68;
        fc1_weights[53][30] = 16'sd26;
        fc1_weights[53][31] = 16'sd17;
        fc1_weights[53][32] = 16'sd14;
        fc1_weights[53][33] = 16'sd43;
        fc1_weights[53][34] = 16'sd35;
        fc1_weights[53][35] = 16'sd-16;
        fc1_weights[53][36] = 16'sd-26;
        fc1_weights[53][37] = 16'sd61;
        fc1_weights[53][38] = 16'sd-47;
        fc1_weights[53][39] = 16'sd-49;
        fc1_weights[53][40] = 16'sd-10;
        fc1_weights[53][41] = 16'sd-63;
        fc1_weights[53][42] = 16'sd45;
        fc1_weights[53][43] = 16'sd10;
        fc1_weights[53][44] = 16'sd-32;
        fc1_weights[53][45] = 16'sd-17;
        fc1_weights[53][46] = 16'sd-21;
        fc1_weights[53][47] = 16'sd-10;
        fc1_weights[53][48] = 16'sd35;
        fc1_weights[53][49] = 16'sd-21;
        fc1_weights[53][50] = 16'sd41;
        fc1_weights[53][51] = 16'sd-7;
        fc1_weights[53][52] = 16'sd25;
        fc1_weights[53][53] = 16'sd-2;
        fc1_weights[53][54] = 16'sd17;
        fc1_weights[53][55] = 16'sd-7;
        fc1_weights[53][56] = 16'sd-2;
        fc1_weights[53][57] = 16'sd-12;
        fc1_weights[53][58] = 16'sd2;
        fc1_weights[53][59] = 16'sd32;
        fc1_weights[53][60] = 16'sd-9;
        fc1_weights[53][61] = 16'sd0;
        fc1_weights[53][62] = 16'sd-24;
        fc1_weights[53][63] = 16'sd18;
        fc1_weights[53][64] = 16'sd-33;
        fc1_weights[53][65] = 16'sd-20;
        fc1_weights[53][66] = 16'sd38;
        fc1_weights[53][67] = 16'sd1;
        fc1_weights[53][68] = 16'sd19;
        fc1_weights[53][69] = 16'sd21;
        fc1_weights[53][70] = 16'sd-36;
        fc1_weights[53][71] = 16'sd9;
        fc1_weights[53][72] = 16'sd-3;
        fc1_weights[53][73] = 16'sd23;
        fc1_weights[53][74] = 16'sd45;
        fc1_weights[53][75] = 16'sd26;
        fc1_weights[53][76] = 16'sd10;
        fc1_weights[53][77] = 16'sd24;
        fc1_weights[53][78] = 16'sd1;
        fc1_weights[53][79] = 16'sd24;
        fc1_weights[53][80] = 16'sd10;
        fc1_weights[53][81] = 16'sd29;
        fc1_weights[53][82] = 16'sd14;
        fc1_weights[53][83] = 16'sd18;
        fc1_weights[53][84] = 16'sd16;
        fc1_weights[53][85] = 16'sd34;
        fc1_weights[53][86] = 16'sd46;
        fc1_weights[53][87] = 16'sd-10;
        fc1_weights[53][88] = 16'sd-2;
        fc1_weights[53][89] = 16'sd14;
        fc1_weights[53][90] = 16'sd-61;
        fc1_weights[53][91] = 16'sd43;
        fc1_weights[53][92] = 16'sd-21;
        fc1_weights[53][93] = 16'sd2;
        fc1_weights[53][94] = 16'sd-17;
        fc1_weights[53][95] = 16'sd-45;
        fc1_weights[53][96] = 16'sd-49;
        fc1_weights[53][97] = 16'sd-39;
        fc1_weights[53][98] = 16'sd-2;
        fc1_weights[53][99] = 16'sd-23;
        fc1_weights[53][100] = 16'sd50;
        fc1_weights[53][101] = 16'sd48;
        fc1_weights[53][102] = 16'sd39;
        fc1_weights[53][103] = 16'sd50;
        fc1_weights[53][104] = 16'sd50;
        fc1_weights[53][105] = 16'sd19;
        fc1_weights[53][106] = 16'sd40;
        fc1_weights[53][107] = 16'sd-39;
        fc1_weights[53][108] = 16'sd2;
        fc1_weights[53][109] = 16'sd-11;
        fc1_weights[53][110] = 16'sd-68;
        fc1_weights[53][111] = 16'sd-21;
        fc1_weights[53][112] = 16'sd-73;
        fc1_weights[53][113] = 16'sd-30;
        fc1_weights[53][114] = 16'sd6;
        fc1_weights[53][115] = 16'sd37;
        fc1_weights[53][116] = 16'sd-56;
        fc1_weights[53][117] = 16'sd-57;
        fc1_weights[53][118] = 16'sd-95;
        fc1_weights[53][119] = 16'sd-66;
        fc1_weights[53][120] = 16'sd-43;
        fc1_weights[53][121] = 16'sd-30;
        fc1_weights[53][122] = 16'sd9;
        fc1_weights[53][123] = 16'sd-26;
        fc1_weights[53][124] = 16'sd-11;
        fc1_weights[53][125] = 16'sd-48;
        fc1_weights[53][126] = 16'sd32;
        fc1_weights[53][127] = 16'sd17;
        fc1_weights[53][128] = 16'sd27;
        fc1_weights[53][129] = 16'sd53;
        fc1_weights[53][130] = 16'sd23;
        fc1_weights[53][131] = 16'sd6;
        fc1_weights[53][132] = 16'sd15;
        fc1_weights[53][133] = 16'sd-10;
        fc1_weights[53][134] = 16'sd19;
        fc1_weights[53][135] = 16'sd-27;
        fc1_weights[53][136] = 16'sd19;
        fc1_weights[53][137] = 16'sd44;
        fc1_weights[53][138] = 16'sd31;
        fc1_weights[53][139] = 16'sd25;
        fc1_weights[53][140] = 16'sd70;
        fc1_weights[53][141] = 16'sd127;
        fc1_weights[53][142] = 16'sd2;
        fc1_weights[53][143] = 16'sd10;
        fc1_weights[53][144] = 16'sd6;
        fc1_weights[53][145] = 16'sd48;
        fc1_weights[53][146] = 16'sd-9;
        fc1_weights[53][147] = 16'sd-24;
        fc1_weights[53][148] = 16'sd-24;
        fc1_weights[53][149] = 16'sd16;
        fc1_weights[53][150] = 16'sd-31;
        fc1_weights[53][151] = 16'sd-28;
        fc1_weights[53][152] = 16'sd-19;
        fc1_weights[53][153] = 16'sd-15;
        fc1_weights[53][154] = 16'sd24;
        fc1_weights[53][155] = 16'sd-22;
        fc1_weights[53][156] = 16'sd42;
        fc1_weights[53][157] = 16'sd-7;
        fc1_weights[53][158] = 16'sd22;
        fc1_weights[53][159] = 16'sd68;
        fc1_weights[53][160] = 16'sd26;
        fc1_weights[53][161] = 16'sd-22;
        fc1_weights[53][162] = 16'sd-20;
        fc1_weights[53][163] = 16'sd-5;
        fc1_weights[53][164] = 16'sd33;
        fc1_weights[53][165] = 16'sd44;
        fc1_weights[53][166] = 16'sd36;
        fc1_weights[53][167] = 16'sd25;
        fc1_weights[53][168] = 16'sd35;
        fc1_weights[53][169] = 16'sd-17;
        fc1_weights[53][170] = 16'sd-51;
        fc1_weights[53][171] = 16'sd-39;
        fc1_weights[53][172] = 16'sd19;
        fc1_weights[53][173] = 16'sd-30;
        fc1_weights[53][174] = 16'sd-23;
        fc1_weights[53][175] = 16'sd-62;
        fc1_weights[53][176] = 16'sd-25;
        fc1_weights[53][177] = 16'sd-23;
        fc1_weights[53][178] = 16'sd11;
        fc1_weights[53][179] = 16'sd20;
        fc1_weights[53][180] = 16'sd27;
        fc1_weights[53][181] = 16'sd51;
        fc1_weights[53][182] = 16'sd24;
        fc1_weights[53][183] = 16'sd20;
        fc1_weights[53][184] = 16'sd-38;
        fc1_weights[53][185] = 16'sd-12;
        fc1_weights[53][186] = 16'sd-4;
        fc1_weights[53][187] = 16'sd-59;
        fc1_weights[53][188] = 16'sd23;
        fc1_weights[53][189] = 16'sd2;
        fc1_weights[53][190] = 16'sd-3;
        fc1_weights[53][191] = 16'sd41;
        fc1_weights[53][192] = 16'sd38;
        fc1_weights[53][193] = 16'sd36;
        fc1_weights[53][194] = 16'sd2;
        fc1_weights[53][195] = 16'sd0;
        fc1_weights[53][196] = 16'sd-32;
        fc1_weights[53][197] = 16'sd-78;
        fc1_weights[53][198] = 16'sd-21;
        fc1_weights[53][199] = 16'sd-32;
        fc1_weights[53][200] = 16'sd-14;
        fc1_weights[53][201] = 16'sd9;
        fc1_weights[53][202] = 16'sd-10;
        fc1_weights[53][203] = 16'sd-21;
        fc1_weights[53][204] = 16'sd-6;
        fc1_weights[53][205] = 16'sd-3;
        fc1_weights[53][206] = 16'sd23;
        fc1_weights[53][207] = 16'sd30;
        fc1_weights[54][0] = 16'sd40;
        fc1_weights[54][1] = 16'sd49;
        fc1_weights[54][2] = 16'sd7;
        fc1_weights[54][3] = 16'sd-38;
        fc1_weights[54][4] = 16'sd-42;
        fc1_weights[54][5] = 16'sd32;
        fc1_weights[54][6] = 16'sd-11;
        fc1_weights[54][7] = 16'sd48;
        fc1_weights[54][8] = 16'sd-90;
        fc1_weights[54][9] = 16'sd-109;
        fc1_weights[54][10] = 16'sd-40;
        fc1_weights[54][11] = 16'sd-46;
        fc1_weights[54][12] = 16'sd15;
        fc1_weights[54][13] = 16'sd67;
        fc1_weights[54][14] = 16'sd66;
        fc1_weights[54][15] = 16'sd14;
        fc1_weights[54][16] = 16'sd40;
        fc1_weights[54][17] = 16'sd43;
        fc1_weights[54][18] = 16'sd-6;
        fc1_weights[54][19] = 16'sd-14;
        fc1_weights[54][20] = 16'sd43;
        fc1_weights[54][21] = 16'sd-16;
        fc1_weights[54][22] = 16'sd20;
        fc1_weights[54][23] = 16'sd49;
        fc1_weights[54][24] = 16'sd65;
        fc1_weights[54][25] = 16'sd61;
        fc1_weights[54][26] = 16'sd24;
        fc1_weights[54][27] = 16'sd6;
        fc1_weights[54][28] = 16'sd-20;
        fc1_weights[54][29] = 16'sd26;
        fc1_weights[54][30] = 16'sd-7;
        fc1_weights[54][31] = 16'sd-25;
        fc1_weights[54][32] = 16'sd1;
        fc1_weights[54][33] = 16'sd-11;
        fc1_weights[54][34] = 16'sd-21;
        fc1_weights[54][35] = 16'sd-27;
        fc1_weights[54][36] = 16'sd-73;
        fc1_weights[54][37] = 16'sd-59;
        fc1_weights[54][38] = 16'sd40;
        fc1_weights[54][39] = 16'sd62;
        fc1_weights[54][40] = 16'sd80;
        fc1_weights[54][41] = 16'sd9;
        fc1_weights[54][42] = 16'sd-67;
        fc1_weights[54][43] = 16'sd-26;
        fc1_weights[54][44] = 16'sd11;
        fc1_weights[54][45] = 16'sd1;
        fc1_weights[54][46] = 16'sd8;
        fc1_weights[54][47] = 16'sd-40;
        fc1_weights[54][48] = 16'sd-63;
        fc1_weights[54][49] = 16'sd21;
        fc1_weights[54][50] = 16'sd21;
        fc1_weights[54][51] = 16'sd45;
        fc1_weights[54][52] = 16'sd-105;
        fc1_weights[54][53] = 16'sd-10;
        fc1_weights[54][54] = 16'sd-47;
        fc1_weights[54][55] = 16'sd-12;
        fc1_weights[54][56] = 16'sd-20;
        fc1_weights[54][57] = 16'sd20;
        fc1_weights[54][58] = 16'sd24;
        fc1_weights[54][59] = 16'sd32;
        fc1_weights[54][60] = 16'sd-14;
        fc1_weights[54][61] = 16'sd-87;
        fc1_weights[54][62] = 16'sd-32;
        fc1_weights[54][63] = 16'sd3;
        fc1_weights[54][64] = 16'sd72;
        fc1_weights[54][65] = 16'sd8;
        fc1_weights[54][66] = 16'sd-5;
        fc1_weights[54][67] = 16'sd-36;
        fc1_weights[54][68] = 16'sd-76;
        fc1_weights[54][69] = 16'sd7;
        fc1_weights[54][70] = 16'sd109;
        fc1_weights[54][71] = 16'sd54;
        fc1_weights[54][72] = 16'sd0;
        fc1_weights[54][73] = 16'sd16;
        fc1_weights[54][74] = 16'sd-23;
        fc1_weights[54][75] = 16'sd-58;
        fc1_weights[54][76] = 16'sd-39;
        fc1_weights[54][77] = 16'sd85;
        fc1_weights[54][78] = 16'sd-71;
        fc1_weights[54][79] = 16'sd5;
        fc1_weights[54][80] = 16'sd-67;
        fc1_weights[54][81] = 16'sd-80;
        fc1_weights[54][82] = 16'sd-51;
        fc1_weights[54][83] = 16'sd28;
        fc1_weights[54][84] = 16'sd-20;
        fc1_weights[54][85] = 16'sd-48;
        fc1_weights[54][86] = 16'sd-46;
        fc1_weights[54][87] = 16'sd9;
        fc1_weights[54][88] = 16'sd15;
        fc1_weights[54][89] = 16'sd-124;
        fc1_weights[54][90] = 16'sd75;
        fc1_weights[54][91] = 16'sd-17;
        fc1_weights[54][92] = 16'sd15;
        fc1_weights[54][93] = 16'sd86;
        fc1_weights[54][94] = 16'sd-22;
        fc1_weights[54][95] = 16'sd-19;
        fc1_weights[54][96] = 16'sd18;
        fc1_weights[54][97] = 16'sd32;
        fc1_weights[54][98] = 16'sd4;
        fc1_weights[54][99] = 16'sd-47;
        fc1_weights[54][100] = 16'sd-43;
        fc1_weights[54][101] = 16'sd-15;
        fc1_weights[54][102] = 16'sd-62;
        fc1_weights[54][103] = 16'sd-38;
        fc1_weights[54][104] = 16'sd-35;
        fc1_weights[54][105] = 16'sd-51;
        fc1_weights[54][106] = 16'sd-13;
        fc1_weights[54][107] = 16'sd-53;
        fc1_weights[54][108] = 16'sd-55;
        fc1_weights[54][109] = 16'sd-15;
        fc1_weights[54][110] = 16'sd-34;
        fc1_weights[54][111] = 16'sd-27;
        fc1_weights[54][112] = 16'sd-7;
        fc1_weights[54][113] = 16'sd-37;
        fc1_weights[54][114] = 16'sd41;
        fc1_weights[54][115] = 16'sd-80;
        fc1_weights[54][116] = 16'sd-33;
        fc1_weights[54][117] = 16'sd-28;
        fc1_weights[54][118] = 16'sd-22;
        fc1_weights[54][119] = 16'sd13;
        fc1_weights[54][120] = 16'sd-1;
        fc1_weights[54][121] = 16'sd-6;
        fc1_weights[54][122] = 16'sd-60;
        fc1_weights[54][123] = 16'sd-7;
        fc1_weights[54][124] = 16'sd-31;
        fc1_weights[54][125] = 16'sd-2;
        fc1_weights[54][126] = 16'sd20;
        fc1_weights[54][127] = 16'sd1;
        fc1_weights[54][128] = 16'sd26;
        fc1_weights[54][129] = 16'sd77;
        fc1_weights[54][130] = 16'sd-49;
        fc1_weights[54][131] = 16'sd46;
        fc1_weights[54][132] = 16'sd38;
        fc1_weights[54][133] = 16'sd59;
        fc1_weights[54][134] = 16'sd88;
        fc1_weights[54][135] = 16'sd51;
        fc1_weights[54][136] = 16'sd45;
        fc1_weights[54][137] = 16'sd-11;
        fc1_weights[54][138] = 16'sd62;
        fc1_weights[54][139] = 16'sd-48;
        fc1_weights[54][140] = 16'sd6;
        fc1_weights[54][141] = 16'sd35;
        fc1_weights[54][142] = 16'sd13;
        fc1_weights[54][143] = 16'sd2;
        fc1_weights[54][144] = 16'sd48;
        fc1_weights[54][145] = 16'sd-18;
        fc1_weights[54][146] = 16'sd-5;
        fc1_weights[54][147] = 16'sd-11;
        fc1_weights[54][148] = 16'sd-12;
        fc1_weights[54][149] = 16'sd21;
        fc1_weights[54][150] = 16'sd43;
        fc1_weights[54][151] = 16'sd105;
        fc1_weights[54][152] = 16'sd-6;
        fc1_weights[54][153] = 16'sd-34;
        fc1_weights[54][154] = 16'sd24;
        fc1_weights[54][155] = 16'sd60;
        fc1_weights[54][156] = 16'sd-28;
        fc1_weights[54][157] = 16'sd28;
        fc1_weights[54][158] = 16'sd19;
        fc1_weights[54][159] = 16'sd46;
        fc1_weights[54][160] = 16'sd13;
        fc1_weights[54][161] = 16'sd64;
        fc1_weights[54][162] = 16'sd74;
        fc1_weights[54][163] = 16'sd46;
        fc1_weights[54][164] = 16'sd29;
        fc1_weights[54][165] = 16'sd-27;
        fc1_weights[54][166] = 16'sd-20;
        fc1_weights[54][167] = 16'sd-18;
        fc1_weights[54][168] = 16'sd-26;
        fc1_weights[54][169] = 16'sd38;
        fc1_weights[54][170] = 16'sd45;
        fc1_weights[54][171] = 16'sd-22;
        fc1_weights[54][172] = 16'sd-7;
        fc1_weights[54][173] = 16'sd-15;
        fc1_weights[54][174] = 16'sd10;
        fc1_weights[54][175] = 16'sd-21;
        fc1_weights[54][176] = 16'sd14;
        fc1_weights[54][177] = 16'sd43;
        fc1_weights[54][178] = 16'sd-16;
        fc1_weights[54][179] = 16'sd38;
        fc1_weights[54][180] = 16'sd2;
        fc1_weights[54][181] = 16'sd-12;
        fc1_weights[54][182] = 16'sd79;
        fc1_weights[54][183] = 16'sd5;
        fc1_weights[54][184] = 16'sd52;
        fc1_weights[54][185] = 16'sd10;
        fc1_weights[54][186] = 16'sd52;
        fc1_weights[54][187] = 16'sd-47;
        fc1_weights[54][188] = 16'sd-17;
        fc1_weights[54][189] = 16'sd7;
        fc1_weights[54][190] = 16'sd41;
        fc1_weights[54][191] = 16'sd-52;
        fc1_weights[54][192] = 16'sd-44;
        fc1_weights[54][193] = 16'sd-16;
        fc1_weights[54][194] = 16'sd-21;
        fc1_weights[54][195] = 16'sd24;
        fc1_weights[54][196] = 16'sd45;
        fc1_weights[54][197] = 16'sd68;
        fc1_weights[54][198] = 16'sd-39;
        fc1_weights[54][199] = 16'sd-52;
        fc1_weights[54][200] = 16'sd48;
        fc1_weights[54][201] = 16'sd-66;
        fc1_weights[54][202] = 16'sd-57;
        fc1_weights[54][203] = 16'sd70;
        fc1_weights[54][204] = 16'sd5;
        fc1_weights[54][205] = 16'sd-5;
        fc1_weights[54][206] = 16'sd-22;
        fc1_weights[54][207] = 16'sd14;
        fc1_weights[55][0] = 16'sd-22;
        fc1_weights[55][1] = 16'sd15;
        fc1_weights[55][2] = 16'sd1;
        fc1_weights[55][3] = 16'sd3;
        fc1_weights[55][4] = 16'sd9;
        fc1_weights[55][5] = 16'sd38;
        fc1_weights[55][6] = 16'sd50;
        fc1_weights[55][7] = 16'sd64;
        fc1_weights[55][8] = 16'sd4;
        fc1_weights[55][9] = 16'sd-76;
        fc1_weights[55][10] = 16'sd-74;
        fc1_weights[55][11] = 16'sd-55;
        fc1_weights[55][12] = 16'sd9;
        fc1_weights[55][13] = 16'sd57;
        fc1_weights[55][14] = 16'sd-18;
        fc1_weights[55][15] = 16'sd-10;
        fc1_weights[55][16] = 16'sd2;
        fc1_weights[55][17] = 16'sd36;
        fc1_weights[55][18] = 16'sd25;
        fc1_weights[55][19] = 16'sd-4;
        fc1_weights[55][20] = 16'sd46;
        fc1_weights[55][21] = 16'sd-19;
        fc1_weights[55][22] = 16'sd10;
        fc1_weights[55][23] = 16'sd23;
        fc1_weights[55][24] = 16'sd9;
        fc1_weights[55][25] = 16'sd42;
        fc1_weights[55][26] = 16'sd27;
        fc1_weights[55][27] = 16'sd-12;
        fc1_weights[55][28] = 16'sd-5;
        fc1_weights[55][29] = 16'sd48;
        fc1_weights[55][30] = 16'sd50;
        fc1_weights[55][31] = 16'sd-3;
        fc1_weights[55][32] = 16'sd16;
        fc1_weights[55][33] = 16'sd-9;
        fc1_weights[55][34] = 16'sd35;
        fc1_weights[55][35] = 16'sd0;
        fc1_weights[55][36] = 16'sd-70;
        fc1_weights[55][37] = 16'sd-39;
        fc1_weights[55][38] = 16'sd-6;
        fc1_weights[55][39] = 16'sd6;
        fc1_weights[55][40] = 16'sd-40;
        fc1_weights[55][41] = 16'sd7;
        fc1_weights[55][42] = 16'sd14;
        fc1_weights[55][43] = 16'sd-13;
        fc1_weights[55][44] = 16'sd-7;
        fc1_weights[55][45] = 16'sd-15;
        fc1_weights[55][46] = 16'sd56;
        fc1_weights[55][47] = 16'sd-21;
        fc1_weights[55][48] = 16'sd2;
        fc1_weights[55][49] = 16'sd6;
        fc1_weights[55][50] = 16'sd8;
        fc1_weights[55][51] = 16'sd19;
        fc1_weights[55][52] = 16'sd-11;
        fc1_weights[55][53] = 16'sd15;
        fc1_weights[55][54] = 16'sd-54;
        fc1_weights[55][55] = 16'sd21;
        fc1_weights[55][56] = 16'sd-12;
        fc1_weights[55][57] = 16'sd12;
        fc1_weights[55][58] = 16'sd-4;
        fc1_weights[55][59] = 16'sd6;
        fc1_weights[55][60] = 16'sd5;
        fc1_weights[55][61] = 16'sd-29;
        fc1_weights[55][62] = 16'sd-60;
        fc1_weights[55][63] = 16'sd-37;
        fc1_weights[55][64] = 16'sd37;
        fc1_weights[55][65] = 16'sd-59;
        fc1_weights[55][66] = 16'sd17;
        fc1_weights[55][67] = 16'sd13;
        fc1_weights[55][68] = 16'sd-14;
        fc1_weights[55][69] = 16'sd37;
        fc1_weights[55][70] = 16'sd41;
        fc1_weights[55][71] = 16'sd24;
        fc1_weights[55][72] = 16'sd14;
        fc1_weights[55][73] = 16'sd56;
        fc1_weights[55][74] = 16'sd26;
        fc1_weights[55][75] = 16'sd5;
        fc1_weights[55][76] = 16'sd-24;
        fc1_weights[55][77] = 16'sd9;
        fc1_weights[55][78] = 16'sd19;
        fc1_weights[55][79] = 16'sd20;
        fc1_weights[55][80] = 16'sd-14;
        fc1_weights[55][81] = 16'sd23;
        fc1_weights[55][82] = 16'sd17;
        fc1_weights[55][83] = 16'sd13;
        fc1_weights[55][84] = 16'sd-25;
        fc1_weights[55][85] = 16'sd-48;
        fc1_weights[55][86] = 16'sd-39;
        fc1_weights[55][87] = 16'sd-45;
        fc1_weights[55][88] = 16'sd-32;
        fc1_weights[55][89] = 16'sd-52;
        fc1_weights[55][90] = 16'sd-40;
        fc1_weights[55][91] = 16'sd-17;
        fc1_weights[55][92] = 16'sd1;
        fc1_weights[55][93] = 16'sd0;
        fc1_weights[55][94] = 16'sd-39;
        fc1_weights[55][95] = 16'sd18;
        fc1_weights[55][96] = 16'sd22;
        fc1_weights[55][97] = 16'sd-4;
        fc1_weights[55][98] = 16'sd27;
        fc1_weights[55][99] = 16'sd5;
        fc1_weights[55][100] = 16'sd23;
        fc1_weights[55][101] = 16'sd16;
        fc1_weights[55][102] = 16'sd-24;
        fc1_weights[55][103] = 16'sd22;
        fc1_weights[55][104] = 16'sd38;
        fc1_weights[55][105] = 16'sd1;
        fc1_weights[55][106] = 16'sd1;
        fc1_weights[55][107] = 16'sd17;
        fc1_weights[55][108] = 16'sd15;
        fc1_weights[55][109] = 16'sd29;
        fc1_weights[55][110] = 16'sd-1;
        fc1_weights[55][111] = 16'sd-16;
        fc1_weights[55][112] = 16'sd-39;
        fc1_weights[55][113] = 16'sd-76;
        fc1_weights[55][114] = 16'sd-24;
        fc1_weights[55][115] = 16'sd-25;
        fc1_weights[55][116] = 16'sd-6;
        fc1_weights[55][117] = 16'sd-8;
        fc1_weights[55][118] = 16'sd7;
        fc1_weights[55][119] = 16'sd-18;
        fc1_weights[55][120] = 16'sd-16;
        fc1_weights[55][121] = 16'sd5;
        fc1_weights[55][122] = 16'sd-45;
        fc1_weights[55][123] = 16'sd-2;
        fc1_weights[55][124] = 16'sd-18;
        fc1_weights[55][125] = 16'sd3;
        fc1_weights[55][126] = 16'sd45;
        fc1_weights[55][127] = 16'sd-6;
        fc1_weights[55][128] = 16'sd24;
        fc1_weights[55][129] = 16'sd62;
        fc1_weights[55][130] = 16'sd12;
        fc1_weights[55][131] = 16'sd18;
        fc1_weights[55][132] = 16'sd-16;
        fc1_weights[55][133] = 16'sd6;
        fc1_weights[55][134] = 16'sd-8;
        fc1_weights[55][135] = 16'sd2;
        fc1_weights[55][136] = 16'sd-7;
        fc1_weights[55][137] = 16'sd-44;
        fc1_weights[55][138] = 16'sd2;
        fc1_weights[55][139] = 16'sd-65;
        fc1_weights[55][140] = 16'sd-11;
        fc1_weights[55][141] = 16'sd35;
        fc1_weights[55][142] = 16'sd-20;
        fc1_weights[55][143] = 16'sd22;
        fc1_weights[55][144] = 16'sd74;
        fc1_weights[55][145] = 16'sd55;
        fc1_weights[55][146] = 16'sd30;
        fc1_weights[55][147] = 16'sd26;
        fc1_weights[55][148] = 16'sd45;
        fc1_weights[55][149] = 16'sd8;
        fc1_weights[55][150] = 16'sd-15;
        fc1_weights[55][151] = 16'sd30;
        fc1_weights[55][152] = 16'sd-13;
        fc1_weights[55][153] = 16'sd-36;
        fc1_weights[55][154] = 16'sd27;
        fc1_weights[55][155] = 16'sd1;
        fc1_weights[55][156] = 16'sd-34;
        fc1_weights[55][157] = 16'sd-1;
        fc1_weights[55][158] = 16'sd-30;
        fc1_weights[55][159] = 16'sd16;
        fc1_weights[55][160] = 16'sd0;
        fc1_weights[55][161] = 16'sd24;
        fc1_weights[55][162] = 16'sd5;
        fc1_weights[55][163] = 16'sd13;
        fc1_weights[55][164] = 16'sd-4;
        fc1_weights[55][165] = 16'sd-46;
        fc1_weights[55][166] = 16'sd-63;
        fc1_weights[55][167] = 16'sd-24;
        fc1_weights[55][168] = 16'sd6;
        fc1_weights[55][169] = 16'sd20;
        fc1_weights[55][170] = 16'sd55;
        fc1_weights[55][171] = 16'sd17;
        fc1_weights[55][172] = 16'sd3;
        fc1_weights[55][173] = 16'sd-1;
        fc1_weights[55][174] = 16'sd20;
        fc1_weights[55][175] = 16'sd-1;
        fc1_weights[55][176] = 16'sd-17;
        fc1_weights[55][177] = 16'sd-9;
        fc1_weights[55][178] = 16'sd19;
        fc1_weights[55][179] = 16'sd-21;
        fc1_weights[55][180] = 16'sd57;
        fc1_weights[55][181] = 16'sd27;
        fc1_weights[55][182] = 16'sd-20;
        fc1_weights[55][183] = 16'sd16;
        fc1_weights[55][184] = 16'sd12;
        fc1_weights[55][185] = 16'sd-16;
        fc1_weights[55][186] = 16'sd-21;
        fc1_weights[55][187] = 16'sd-47;
        fc1_weights[55][188] = 16'sd-53;
        fc1_weights[55][189] = 16'sd-6;
        fc1_weights[55][190] = 16'sd-2;
        fc1_weights[55][191] = 16'sd-17;
        fc1_weights[55][192] = 16'sd16;
        fc1_weights[55][193] = 16'sd8;
        fc1_weights[55][194] = 16'sd10;
        fc1_weights[55][195] = 16'sd25;
        fc1_weights[55][196] = 16'sd37;
        fc1_weights[55][197] = 16'sd7;
        fc1_weights[55][198] = 16'sd7;
        fc1_weights[55][199] = 16'sd-12;
        fc1_weights[55][200] = 16'sd7;
        fc1_weights[55][201] = 16'sd-4;
        fc1_weights[55][202] = 16'sd15;
        fc1_weights[55][203] = 16'sd-21;
        fc1_weights[55][204] = 16'sd-11;
        fc1_weights[55][205] = 16'sd-3;
        fc1_weights[55][206] = 16'sd-1;
        fc1_weights[55][207] = 16'sd58;
        fc1_weights[56][0] = 16'sd-23;
        fc1_weights[56][1] = 16'sd-13;
        fc1_weights[56][2] = 16'sd-35;
        fc1_weights[56][3] = 16'sd-28;
        fc1_weights[56][4] = 16'sd-31;
        fc1_weights[56][5] = 16'sd-26;
        fc1_weights[56][6] = 16'sd-50;
        fc1_weights[56][7] = 16'sd-39;
        fc1_weights[56][8] = 16'sd-40;
        fc1_weights[56][9] = 16'sd-51;
        fc1_weights[56][10] = 16'sd-1;
        fc1_weights[56][11] = 16'sd-46;
        fc1_weights[56][12] = 16'sd-19;
        fc1_weights[56][13] = 16'sd-3;
        fc1_weights[56][14] = 16'sd-3;
        fc1_weights[56][15] = 16'sd38;
        fc1_weights[56][16] = 16'sd27;
        fc1_weights[56][17] = 16'sd-18;
        fc1_weights[56][18] = 16'sd4;
        fc1_weights[56][19] = 16'sd-14;
        fc1_weights[56][20] = 16'sd13;
        fc1_weights[56][21] = 16'sd-29;
        fc1_weights[56][22] = 16'sd-9;
        fc1_weights[56][23] = 16'sd-15;
        fc1_weights[56][24] = 16'sd0;
        fc1_weights[56][25] = 16'sd3;
        fc1_weights[56][26] = 16'sd-9;
        fc1_weights[56][27] = 16'sd-11;
        fc1_weights[56][28] = 16'sd-3;
        fc1_weights[56][29] = 16'sd1;
        fc1_weights[56][30] = 16'sd6;
        fc1_weights[56][31] = 16'sd10;
        fc1_weights[56][32] = 16'sd-24;
        fc1_weights[56][33] = 16'sd-48;
        fc1_weights[56][34] = 16'sd-53;
        fc1_weights[56][35] = 16'sd-54;
        fc1_weights[56][36] = 16'sd-34;
        fc1_weights[56][37] = 16'sd-53;
        fc1_weights[56][38] = 16'sd-48;
        fc1_weights[56][39] = 16'sd1;
        fc1_weights[56][40] = 16'sd9;
        fc1_weights[56][41] = 16'sd55;
        fc1_weights[56][42] = 16'sd-6;
        fc1_weights[56][43] = 16'sd-27;
        fc1_weights[56][44] = 16'sd1;
        fc1_weights[56][45] = 16'sd-36;
        fc1_weights[56][46] = 16'sd-27;
        fc1_weights[56][47] = 16'sd1;
        fc1_weights[56][48] = 16'sd-2;
        fc1_weights[56][49] = 16'sd4;
        fc1_weights[56][50] = 16'sd14;
        fc1_weights[56][51] = 16'sd-17;
        fc1_weights[56][52] = 16'sd7;
        fc1_weights[56][53] = 16'sd19;
        fc1_weights[56][54] = 16'sd12;
        fc1_weights[56][55] = 16'sd-17;
        fc1_weights[56][56] = 16'sd42;
        fc1_weights[56][57] = 16'sd20;
        fc1_weights[56][58] = 16'sd7;
        fc1_weights[56][59] = 16'sd7;
        fc1_weights[56][60] = 16'sd6;
        fc1_weights[56][61] = 16'sd-1;
        fc1_weights[56][62] = 16'sd-42;
        fc1_weights[56][63] = 16'sd-53;
        fc1_weights[56][64] = 16'sd-35;
        fc1_weights[56][65] = 16'sd-5;
        fc1_weights[56][66] = 16'sd24;
        fc1_weights[56][67] = 16'sd4;
        fc1_weights[56][68] = 16'sd8;
        fc1_weights[56][69] = 16'sd-18;
        fc1_weights[56][70] = 16'sd3;
        fc1_weights[56][71] = 16'sd20;
        fc1_weights[56][72] = 16'sd18;
        fc1_weights[56][73] = 16'sd-13;
        fc1_weights[56][74] = 16'sd0;
        fc1_weights[56][75] = 16'sd-1;
        fc1_weights[56][76] = 16'sd-14;
        fc1_weights[56][77] = 16'sd3;
        fc1_weights[56][78] = 16'sd21;
        fc1_weights[56][79] = 16'sd49;
        fc1_weights[56][80] = 16'sd-6;
        fc1_weights[56][81] = 16'sd18;
        fc1_weights[56][82] = 16'sd9;
        fc1_weights[56][83] = 16'sd3;
        fc1_weights[56][84] = 16'sd2;
        fc1_weights[56][85] = 16'sd0;
        fc1_weights[56][86] = 16'sd4;
        fc1_weights[56][87] = 16'sd10;
        fc1_weights[56][88] = 16'sd3;
        fc1_weights[56][89] = 16'sd-12;
        fc1_weights[56][90] = 16'sd18;
        fc1_weights[56][91] = 16'sd19;
        fc1_weights[56][92] = 16'sd7;
        fc1_weights[56][93] = 16'sd-13;
        fc1_weights[56][94] = 16'sd6;
        fc1_weights[56][95] = 16'sd18;
        fc1_weights[56][96] = 16'sd-4;
        fc1_weights[56][97] = 16'sd-16;
        fc1_weights[56][98] = 16'sd8;
        fc1_weights[56][99] = 16'sd4;
        fc1_weights[56][100] = 16'sd13;
        fc1_weights[56][101] = 16'sd18;
        fc1_weights[56][102] = 16'sd11;
        fc1_weights[56][103] = 16'sd-16;
        fc1_weights[56][104] = 16'sd28;
        fc1_weights[56][105] = 16'sd-13;
        fc1_weights[56][106] = 16'sd-15;
        fc1_weights[56][107] = 16'sd9;
        fc1_weights[56][108] = 16'sd9;
        fc1_weights[56][109] = 16'sd-1;
        fc1_weights[56][110] = 16'sd-1;
        fc1_weights[56][111] = 16'sd5;
        fc1_weights[56][112] = 16'sd44;
        fc1_weights[56][113] = 16'sd13;
        fc1_weights[56][114] = 16'sd-17;
        fc1_weights[56][115] = 16'sd16;
        fc1_weights[56][116] = 16'sd-11;
        fc1_weights[56][117] = 16'sd-18;
        fc1_weights[56][118] = 16'sd22;
        fc1_weights[56][119] = 16'sd21;
        fc1_weights[56][120] = 16'sd27;
        fc1_weights[56][121] = 16'sd-12;
        fc1_weights[56][122] = 16'sd4;
        fc1_weights[56][123] = 16'sd-6;
        fc1_weights[56][124] = 16'sd-32;
        fc1_weights[56][125] = 16'sd-22;
        fc1_weights[56][126] = 16'sd-34;
        fc1_weights[56][127] = 16'sd6;
        fc1_weights[56][128] = 16'sd-14;
        fc1_weights[56][129] = 16'sd-61;
        fc1_weights[56][130] = 16'sd3;
        fc1_weights[56][131] = 16'sd-21;
        fc1_weights[56][132] = 16'sd-1;
        fc1_weights[56][133] = 16'sd15;
        fc1_weights[56][134] = 16'sd13;
        fc1_weights[56][135] = 16'sd-29;
        fc1_weights[56][136] = 16'sd-11;
        fc1_weights[56][137] = 16'sd11;
        fc1_weights[56][138] = 16'sd-27;
        fc1_weights[56][139] = 16'sd2;
        fc1_weights[56][140] = 16'sd-22;
        fc1_weights[56][141] = 16'sd-5;
        fc1_weights[56][142] = 16'sd34;
        fc1_weights[56][143] = 16'sd-17;
        fc1_weights[56][144] = 16'sd-21;
        fc1_weights[56][145] = 16'sd-23;
        fc1_weights[56][146] = 16'sd-24;
        fc1_weights[56][147] = 16'sd9;
        fc1_weights[56][148] = 16'sd-18;
        fc1_weights[56][149] = 16'sd-26;
        fc1_weights[56][150] = 16'sd-23;
        fc1_weights[56][151] = 16'sd14;
        fc1_weights[56][152] = 16'sd7;
        fc1_weights[56][153] = 16'sd27;
        fc1_weights[56][154] = 16'sd-4;
        fc1_weights[56][155] = 16'sd-1;
        fc1_weights[56][156] = 16'sd-16;
        fc1_weights[56][157] = 16'sd-17;
        fc1_weights[56][158] = 16'sd-13;
        fc1_weights[56][159] = 16'sd4;
        fc1_weights[56][160] = 16'sd-18;
        fc1_weights[56][161] = 16'sd-20;
        fc1_weights[56][162] = 16'sd16;
        fc1_weights[56][163] = 16'sd-23;
        fc1_weights[56][164] = 16'sd-36;
        fc1_weights[56][165] = 16'sd-26;
        fc1_weights[56][166] = 16'sd-4;
        fc1_weights[56][167] = 16'sd6;
        fc1_weights[56][168] = 16'sd1;
        fc1_weights[56][169] = 16'sd11;
        fc1_weights[56][170] = 16'sd8;
        fc1_weights[56][171] = 16'sd1;
        fc1_weights[56][172] = 16'sd-29;
        fc1_weights[56][173] = 16'sd-3;
        fc1_weights[56][174] = 16'sd-22;
        fc1_weights[56][175] = 16'sd-6;
        fc1_weights[56][176] = 16'sd-15;
        fc1_weights[56][177] = 16'sd-11;
        fc1_weights[56][178] = 16'sd-26;
        fc1_weights[56][179] = 16'sd-14;
        fc1_weights[56][180] = 16'sd-19;
        fc1_weights[56][181] = 16'sd-11;
        fc1_weights[56][182] = 16'sd4;
        fc1_weights[56][183] = 16'sd-21;
        fc1_weights[56][184] = 16'sd5;
        fc1_weights[56][185] = 16'sd-3;
        fc1_weights[56][186] = 16'sd-32;
        fc1_weights[56][187] = 16'sd-18;
        fc1_weights[56][188] = 16'sd-52;
        fc1_weights[56][189] = 16'sd-20;
        fc1_weights[56][190] = 16'sd5;
        fc1_weights[56][191] = 16'sd12;
        fc1_weights[56][192] = 16'sd13;
        fc1_weights[56][193] = 16'sd26;
        fc1_weights[56][194] = 16'sd44;
        fc1_weights[56][195] = 16'sd24;
        fc1_weights[56][196] = 16'sd14;
        fc1_weights[56][197] = 16'sd15;
        fc1_weights[56][198] = 16'sd7;
        fc1_weights[56][199] = 16'sd48;
        fc1_weights[56][200] = 16'sd8;
        fc1_weights[56][201] = 16'sd-12;
        fc1_weights[56][202] = 16'sd-18;
        fc1_weights[56][203] = 16'sd13;
        fc1_weights[56][204] = 16'sd-8;
        fc1_weights[56][205] = 16'sd-17;
        fc1_weights[56][206] = 16'sd-35;
        fc1_weights[56][207] = 16'sd-1;
        fc1_weights[57][0] = 16'sd-23;
        fc1_weights[57][1] = 16'sd-50;
        fc1_weights[57][2] = 16'sd-46;
        fc1_weights[57][3] = 16'sd-15;
        fc1_weights[57][4] = 16'sd-40;
        fc1_weights[57][5] = 16'sd-36;
        fc1_weights[57][6] = 16'sd15;
        fc1_weights[57][7] = 16'sd22;
        fc1_weights[57][8] = 16'sd14;
        fc1_weights[57][9] = 16'sd15;
        fc1_weights[57][10] = 16'sd20;
        fc1_weights[57][11] = 16'sd46;
        fc1_weights[57][12] = 16'sd-63;
        fc1_weights[57][13] = 16'sd-62;
        fc1_weights[57][14] = 16'sd-7;
        fc1_weights[57][15] = 16'sd72;
        fc1_weights[57][16] = 16'sd75;
        fc1_weights[57][17] = 16'sd-1;
        fc1_weights[57][18] = 16'sd18;
        fc1_weights[57][19] = 16'sd-32;
        fc1_weights[57][20] = 16'sd13;
        fc1_weights[57][21] = 16'sd-67;
        fc1_weights[57][22] = 16'sd-42;
        fc1_weights[57][23] = 16'sd-55;
        fc1_weights[57][24] = 16'sd30;
        fc1_weights[57][25] = 16'sd33;
        fc1_weights[57][26] = 16'sd-54;
        fc1_weights[57][27] = 16'sd-61;
        fc1_weights[57][28] = 16'sd-87;
        fc1_weights[57][29] = 16'sd-9;
        fc1_weights[57][30] = 16'sd45;
        fc1_weights[57][31] = 16'sd3;
        fc1_weights[57][32] = 16'sd-36;
        fc1_weights[57][33] = 16'sd-28;
        fc1_weights[57][34] = 16'sd35;
        fc1_weights[57][35] = 16'sd-11;
        fc1_weights[57][36] = 16'sd40;
        fc1_weights[57][37] = 16'sd37;
        fc1_weights[57][38] = 16'sd-6;
        fc1_weights[57][39] = 16'sd-123;
        fc1_weights[57][40] = 16'sd77;
        fc1_weights[57][41] = 16'sd84;
        fc1_weights[57][42] = 16'sd5;
        fc1_weights[57][43] = 16'sd26;
        fc1_weights[57][44] = 16'sd-4;
        fc1_weights[57][45] = 16'sd-67;
        fc1_weights[57][46] = 16'sd-31;
        fc1_weights[57][47] = 16'sd-39;
        fc1_weights[57][48] = 16'sd0;
        fc1_weights[57][49] = 16'sd15;
        fc1_weights[57][50] = 16'sd0;
        fc1_weights[57][51] = 16'sd-31;
        fc1_weights[57][52] = 16'sd-80;
        fc1_weights[57][53] = 16'sd-20;
        fc1_weights[57][54] = 16'sd33;
        fc1_weights[57][55] = 16'sd28;
        fc1_weights[57][56] = 16'sd-10;
        fc1_weights[57][57] = 16'sd-14;
        fc1_weights[57][58] = 16'sd-7;
        fc1_weights[57][59] = 16'sd-55;
        fc1_weights[57][60] = 16'sd41;
        fc1_weights[57][61] = 16'sd1;
        fc1_weights[57][62] = 16'sd-9;
        fc1_weights[57][63] = 16'sd2;
        fc1_weights[57][64] = 16'sd0;
        fc1_weights[57][65] = 16'sd48;
        fc1_weights[57][66] = 16'sd73;
        fc1_weights[57][67] = 16'sd11;
        fc1_weights[57][68] = 16'sd-3;
        fc1_weights[57][69] = 16'sd-38;
        fc1_weights[57][70] = 16'sd-45;
        fc1_weights[57][71] = 16'sd-23;
        fc1_weights[57][72] = 16'sd20;
        fc1_weights[57][73] = 16'sd-102;
        fc1_weights[57][74] = 16'sd-33;
        fc1_weights[57][75] = 16'sd-22;
        fc1_weights[57][76] = 16'sd38;
        fc1_weights[57][77] = 16'sd53;
        fc1_weights[57][78] = 16'sd-28;
        fc1_weights[57][79] = 16'sd48;
        fc1_weights[57][80] = 16'sd23;
        fc1_weights[57][81] = 16'sd5;
        fc1_weights[57][82] = 16'sd-37;
        fc1_weights[57][83] = 16'sd-44;
        fc1_weights[57][84] = 16'sd-5;
        fc1_weights[57][85] = 16'sd-36;
        fc1_weights[57][86] = 16'sd-20;
        fc1_weights[57][87] = 16'sd16;
        fc1_weights[57][88] = 16'sd-42;
        fc1_weights[57][89] = 16'sd73;
        fc1_weights[57][90] = 16'sd21;
        fc1_weights[57][91] = 16'sd39;
        fc1_weights[57][92] = 16'sd-27;
        fc1_weights[57][93] = 16'sd32;
        fc1_weights[57][94] = 16'sd8;
        fc1_weights[57][95] = 16'sd-9;
        fc1_weights[57][96] = 16'sd-9;
        fc1_weights[57][97] = 16'sd23;
        fc1_weights[57][98] = 16'sd-27;
        fc1_weights[57][99] = 16'sd-5;
        fc1_weights[57][100] = 16'sd-1;
        fc1_weights[57][101] = 16'sd18;
        fc1_weights[57][102] = 16'sd50;
        fc1_weights[57][103] = 16'sd34;
        fc1_weights[57][104] = 16'sd-48;
        fc1_weights[57][105] = 16'sd13;
        fc1_weights[57][106] = 16'sd-18;
        fc1_weights[57][107] = 16'sd-71;
        fc1_weights[57][108] = 16'sd19;
        fc1_weights[57][109] = 16'sd12;
        fc1_weights[57][110] = 16'sd16;
        fc1_weights[57][111] = 16'sd-52;
        fc1_weights[57][112] = 16'sd22;
        fc1_weights[57][113] = 16'sd80;
        fc1_weights[57][114] = 16'sd6;
        fc1_weights[57][115] = 16'sd21;
        fc1_weights[57][116] = 16'sd24;
        fc1_weights[57][117] = 16'sd77;
        fc1_weights[57][118] = 16'sd34;
        fc1_weights[57][119] = 16'sd18;
        fc1_weights[57][120] = 16'sd37;
        fc1_weights[57][121] = 16'sd28;
        fc1_weights[57][122] = 16'sd31;
        fc1_weights[57][123] = 16'sd65;
        fc1_weights[57][124] = 16'sd-47;
        fc1_weights[57][125] = 16'sd-4;
        fc1_weights[57][126] = 16'sd-17;
        fc1_weights[57][127] = 16'sd7;
        fc1_weights[57][128] = 16'sd0;
        fc1_weights[57][129] = 16'sd-66;
        fc1_weights[57][130] = 16'sd-56;
        fc1_weights[57][131] = 16'sd-78;
        fc1_weights[57][132] = 16'sd-15;
        fc1_weights[57][133] = 16'sd-32;
        fc1_weights[57][134] = 16'sd3;
        fc1_weights[57][135] = 16'sd14;
        fc1_weights[57][136] = 16'sd-53;
        fc1_weights[57][137] = 16'sd-52;
        fc1_weights[57][138] = 16'sd24;
        fc1_weights[57][139] = 16'sd42;
        fc1_weights[57][140] = 16'sd67;
        fc1_weights[57][141] = 16'sd-43;
        fc1_weights[57][142] = 16'sd98;
        fc1_weights[57][143] = 16'sd44;
        fc1_weights[57][144] = 16'sd73;
        fc1_weights[57][145] = 16'sd13;
        fc1_weights[57][146] = 16'sd-24;
        fc1_weights[57][147] = 16'sd-22;
        fc1_weights[57][148] = 16'sd4;
        fc1_weights[57][149] = 16'sd-12;
        fc1_weights[57][150] = 16'sd-28;
        fc1_weights[57][151] = 16'sd-14;
        fc1_weights[57][152] = 16'sd11;
        fc1_weights[57][153] = 16'sd25;
        fc1_weights[57][154] = 16'sd4;
        fc1_weights[57][155] = 16'sd19;
        fc1_weights[57][156] = 16'sd32;
        fc1_weights[57][157] = 16'sd-11;
        fc1_weights[57][158] = 16'sd1;
        fc1_weights[57][159] = 16'sd-78;
        fc1_weights[57][160] = 16'sd-74;
        fc1_weights[57][161] = 16'sd-101;
        fc1_weights[57][162] = 16'sd11;
        fc1_weights[57][163] = 16'sd6;
        fc1_weights[57][164] = 16'sd21;
        fc1_weights[57][165] = 16'sd92;
        fc1_weights[57][166] = 16'sd36;
        fc1_weights[57][167] = 16'sd50;
        fc1_weights[57][168] = 16'sd112;
        fc1_weights[57][169] = 16'sd5;
        fc1_weights[57][170] = 16'sd24;
        fc1_weights[57][171] = 16'sd-6;
        fc1_weights[57][172] = 16'sd29;
        fc1_weights[57][173] = 16'sd21;
        fc1_weights[57][174] = 16'sd14;
        fc1_weights[57][175] = 16'sd41;
        fc1_weights[57][176] = 16'sd11;
        fc1_weights[57][177] = 16'sd11;
        fc1_weights[57][178] = 16'sd-35;
        fc1_weights[57][179] = 16'sd45;
        fc1_weights[57][180] = 16'sd36;
        fc1_weights[57][181] = 16'sd45;
        fc1_weights[57][182] = 16'sd-33;
        fc1_weights[57][183] = 16'sd-13;
        fc1_weights[57][184] = 16'sd-50;
        fc1_weights[57][185] = 16'sd-42;
        fc1_weights[57][186] = 16'sd-36;
        fc1_weights[57][187] = 16'sd-10;
        fc1_weights[57][188] = 16'sd33;
        fc1_weights[57][189] = 16'sd-63;
        fc1_weights[57][190] = 16'sd25;
        fc1_weights[57][191] = 16'sd52;
        fc1_weights[57][192] = 16'sd-36;
        fc1_weights[57][193] = 16'sd17;
        fc1_weights[57][194] = 16'sd-16;
        fc1_weights[57][195] = 16'sd26;
        fc1_weights[57][196] = 16'sd-33;
        fc1_weights[57][197] = 16'sd44;
        fc1_weights[57][198] = 16'sd28;
        fc1_weights[57][199] = 16'sd39;
        fc1_weights[57][200] = 16'sd-19;
        fc1_weights[57][201] = 16'sd16;
        fc1_weights[57][202] = 16'sd-24;
        fc1_weights[57][203] = 16'sd48;
        fc1_weights[57][204] = 16'sd16;
        fc1_weights[57][205] = 16'sd2;
        fc1_weights[57][206] = 16'sd-37;
        fc1_weights[57][207] = 16'sd-43;
        fc1_weights[58][0] = 16'sd4;
        fc1_weights[58][1] = 16'sd-17;
        fc1_weights[58][2] = 16'sd-23;
        fc1_weights[58][3] = 16'sd-32;
        fc1_weights[58][4] = 16'sd-16;
        fc1_weights[58][5] = 16'sd-32;
        fc1_weights[58][6] = 16'sd-2;
        fc1_weights[58][7] = 16'sd-35;
        fc1_weights[58][8] = 16'sd-37;
        fc1_weights[58][9] = 16'sd-7;
        fc1_weights[58][10] = 16'sd-32;
        fc1_weights[58][11] = 16'sd-35;
        fc1_weights[58][12] = 16'sd-61;
        fc1_weights[58][13] = 16'sd-37;
        fc1_weights[58][14] = 16'sd9;
        fc1_weights[58][15] = 16'sd8;
        fc1_weights[58][16] = 16'sd21;
        fc1_weights[58][17] = 16'sd-25;
        fc1_weights[58][18] = 16'sd0;
        fc1_weights[58][19] = 16'sd-21;
        fc1_weights[58][20] = 16'sd25;
        fc1_weights[58][21] = 16'sd37;
        fc1_weights[58][22] = 16'sd26;
        fc1_weights[58][23] = 16'sd4;
        fc1_weights[58][24] = 16'sd-2;
        fc1_weights[58][25] = 16'sd22;
        fc1_weights[58][26] = 16'sd-3;
        fc1_weights[58][27] = 16'sd-9;
        fc1_weights[58][28] = 16'sd-6;
        fc1_weights[58][29] = 16'sd-32;
        fc1_weights[58][30] = 16'sd7;
        fc1_weights[58][31] = 16'sd-5;
        fc1_weights[58][32] = 16'sd-30;
        fc1_weights[58][33] = 16'sd-11;
        fc1_weights[58][34] = 16'sd-25;
        fc1_weights[58][35] = 16'sd-19;
        fc1_weights[58][36] = 16'sd-14;
        fc1_weights[58][37] = 16'sd-29;
        fc1_weights[58][38] = 16'sd4;
        fc1_weights[58][39] = 16'sd-11;
        fc1_weights[58][40] = 16'sd27;
        fc1_weights[58][41] = 16'sd12;
        fc1_weights[58][42] = 16'sd-12;
        fc1_weights[58][43] = 16'sd8;
        fc1_weights[58][44] = 16'sd-30;
        fc1_weights[58][45] = 16'sd-51;
        fc1_weights[58][46] = 16'sd-7;
        fc1_weights[58][47] = 16'sd10;
        fc1_weights[58][48] = 16'sd-3;
        fc1_weights[58][49] = 16'sd-12;
        fc1_weights[58][50] = 16'sd-8;
        fc1_weights[58][51] = 16'sd-14;
        fc1_weights[58][52] = 16'sd-7;
        fc1_weights[58][53] = 16'sd-9;
        fc1_weights[58][54] = 16'sd-21;
        fc1_weights[58][55] = 16'sd-32;
        fc1_weights[58][56] = 16'sd-35;
        fc1_weights[58][57] = 16'sd-4;
        fc1_weights[58][58] = 16'sd-1;
        fc1_weights[58][59] = 16'sd-34;
        fc1_weights[58][60] = 16'sd-48;
        fc1_weights[58][61] = 16'sd-37;
        fc1_weights[58][62] = 16'sd-27;
        fc1_weights[58][63] = 16'sd-58;
        fc1_weights[58][64] = 16'sd48;
        fc1_weights[58][65] = 16'sd-46;
        fc1_weights[58][66] = 16'sd11;
        fc1_weights[58][67] = 16'sd2;
        fc1_weights[58][68] = 16'sd-33;
        fc1_weights[58][69] = 16'sd-36;
        fc1_weights[58][70] = 16'sd-57;
        fc1_weights[58][71] = 16'sd17;
        fc1_weights[58][72] = 16'sd42;
        fc1_weights[58][73] = 16'sd-14;
        fc1_weights[58][74] = 16'sd4;
        fc1_weights[58][75] = 16'sd6;
        fc1_weights[58][76] = 16'sd-4;
        fc1_weights[58][77] = 16'sd11;
        fc1_weights[58][78] = 16'sd15;
        fc1_weights[58][79] = 16'sd39;
        fc1_weights[58][80] = 16'sd11;
        fc1_weights[58][81] = 16'sd8;
        fc1_weights[58][82] = 16'sd11;
        fc1_weights[58][83] = 16'sd-13;
        fc1_weights[58][84] = 16'sd28;
        fc1_weights[58][85] = 16'sd-2;
        fc1_weights[58][86] = 16'sd-11;
        fc1_weights[58][87] = 16'sd-32;
        fc1_weights[58][88] = 16'sd-34;
        fc1_weights[58][89] = 16'sd-7;
        fc1_weights[58][90] = 16'sd8;
        fc1_weights[58][91] = 16'sd26;
        fc1_weights[58][92] = 16'sd38;
        fc1_weights[58][93] = 16'sd30;
        fc1_weights[58][94] = 16'sd-18;
        fc1_weights[58][95] = 16'sd16;
        fc1_weights[58][96] = 16'sd-31;
        fc1_weights[58][97] = 16'sd17;
        fc1_weights[58][98] = 16'sd38;
        fc1_weights[58][99] = 16'sd-2;
        fc1_weights[58][100] = 16'sd11;
        fc1_weights[58][101] = 16'sd-31;
        fc1_weights[58][102] = 16'sd-15;
        fc1_weights[58][103] = 16'sd-49;
        fc1_weights[58][104] = 16'sd3;
        fc1_weights[58][105] = 16'sd-16;
        fc1_weights[58][106] = 16'sd15;
        fc1_weights[58][107] = 16'sd-12;
        fc1_weights[58][108] = 16'sd1;
        fc1_weights[58][109] = 16'sd19;
        fc1_weights[58][110] = 16'sd18;
        fc1_weights[58][111] = 16'sd28;
        fc1_weights[58][112] = 16'sd38;
        fc1_weights[58][113] = 16'sd9;
        fc1_weights[58][114] = 16'sd-39;
        fc1_weights[58][115] = 16'sd-48;
        fc1_weights[58][116] = 16'sd-6;
        fc1_weights[58][117] = 16'sd-9;
        fc1_weights[58][118] = 16'sd-4;
        fc1_weights[58][119] = 16'sd10;
        fc1_weights[58][120] = 16'sd-10;
        fc1_weights[58][121] = 16'sd24;
        fc1_weights[58][122] = 16'sd-25;
        fc1_weights[58][123] = 16'sd-10;
        fc1_weights[58][124] = 16'sd11;
        fc1_weights[58][125] = 16'sd-8;
        fc1_weights[58][126] = 16'sd-48;
        fc1_weights[58][127] = 16'sd-11;
        fc1_weights[58][128] = 16'sd14;
        fc1_weights[58][129] = 16'sd-16;
        fc1_weights[58][130] = 16'sd-38;
        fc1_weights[58][131] = 16'sd-45;
        fc1_weights[58][132] = 16'sd-58;
        fc1_weights[58][133] = 16'sd-57;
        fc1_weights[58][134] = 16'sd5;
        fc1_weights[58][135] = 16'sd-1;
        fc1_weights[58][136] = 16'sd29;
        fc1_weights[58][137] = 16'sd13;
        fc1_weights[58][138] = 16'sd14;
        fc1_weights[58][139] = 16'sd82;
        fc1_weights[58][140] = 16'sd58;
        fc1_weights[58][141] = 16'sd13;
        fc1_weights[58][142] = 16'sd16;
        fc1_weights[58][143] = 16'sd-13;
        fc1_weights[58][144] = 16'sd-2;
        fc1_weights[58][145] = 16'sd-5;
        fc1_weights[58][146] = 16'sd-29;
        fc1_weights[58][147] = 16'sd43;
        fc1_weights[58][148] = 16'sd-4;
        fc1_weights[58][149] = 16'sd-20;
        fc1_weights[58][150] = 16'sd-11;
        fc1_weights[58][151] = 16'sd-14;
        fc1_weights[58][152] = 16'sd20;
        fc1_weights[58][153] = 16'sd26;
        fc1_weights[58][154] = 16'sd-5;
        fc1_weights[58][155] = 16'sd10;
        fc1_weights[58][156] = 16'sd18;
        fc1_weights[58][157] = 16'sd26;
        fc1_weights[58][158] = 16'sd12;
        fc1_weights[58][159] = 16'sd9;
        fc1_weights[58][160] = 16'sd33;
        fc1_weights[58][161] = 16'sd21;
        fc1_weights[58][162] = 16'sd-17;
        fc1_weights[58][163] = 16'sd42;
        fc1_weights[58][164] = 16'sd52;
        fc1_weights[58][165] = 16'sd37;
        fc1_weights[58][166] = 16'sd65;
        fc1_weights[58][167] = 16'sd47;
        fc1_weights[58][168] = 16'sd33;
        fc1_weights[58][169] = 16'sd21;
        fc1_weights[58][170] = 16'sd19;
        fc1_weights[58][171] = 16'sd10;
        fc1_weights[58][172] = 16'sd34;
        fc1_weights[58][173] = 16'sd4;
        fc1_weights[58][174] = 16'sd-13;
        fc1_weights[58][175] = 16'sd-17;
        fc1_weights[58][176] = 16'sd-10;
        fc1_weights[58][177] = 16'sd-29;
        fc1_weights[58][178] = 16'sd-36;
        fc1_weights[58][179] = 16'sd-20;
        fc1_weights[58][180] = 16'sd-23;
        fc1_weights[58][181] = 16'sd-15;
        fc1_weights[58][182] = 16'sd-2;
        fc1_weights[58][183] = 16'sd16;
        fc1_weights[58][184] = 16'sd-16;
        fc1_weights[58][185] = 16'sd7;
        fc1_weights[58][186] = 16'sd6;
        fc1_weights[58][187] = 16'sd28;
        fc1_weights[58][188] = 16'sd32;
        fc1_weights[58][189] = 16'sd51;
        fc1_weights[58][190] = 16'sd88;
        fc1_weights[58][191] = 16'sd81;
        fc1_weights[58][192] = 16'sd23;
        fc1_weights[58][193] = 16'sd34;
        fc1_weights[58][194] = 16'sd50;
        fc1_weights[58][195] = 16'sd13;
        fc1_weights[58][196] = 16'sd-21;
        fc1_weights[58][197] = 16'sd-32;
        fc1_weights[58][198] = 16'sd-4;
        fc1_weights[58][199] = 16'sd2;
        fc1_weights[58][200] = 16'sd34;
        fc1_weights[58][201] = 16'sd9;
        fc1_weights[58][202] = 16'sd-33;
        fc1_weights[58][203] = 16'sd27;
        fc1_weights[58][204] = 16'sd0;
        fc1_weights[58][205] = 16'sd13;
        fc1_weights[58][206] = 16'sd36;
        fc1_weights[58][207] = 16'sd-20;
        fc1_weights[59][0] = 16'sd44;
        fc1_weights[59][1] = 16'sd-14;
        fc1_weights[59][2] = 16'sd-55;
        fc1_weights[59][3] = 16'sd22;
        fc1_weights[59][4] = 16'sd-24;
        fc1_weights[59][5] = 16'sd-1;
        fc1_weights[59][6] = 16'sd51;
        fc1_weights[59][7] = 16'sd92;
        fc1_weights[59][8] = 16'sd22;
        fc1_weights[59][9] = 16'sd36;
        fc1_weights[59][10] = 16'sd50;
        fc1_weights[59][11] = 16'sd22;
        fc1_weights[59][12] = 16'sd-32;
        fc1_weights[59][13] = 16'sd-34;
        fc1_weights[59][14] = 16'sd-29;
        fc1_weights[59][15] = 16'sd19;
        fc1_weights[59][16] = 16'sd-7;
        fc1_weights[59][17] = 16'sd-69;
        fc1_weights[59][18] = 16'sd-23;
        fc1_weights[59][19] = 16'sd-33;
        fc1_weights[59][20] = 16'sd-25;
        fc1_weights[59][21] = 16'sd-19;
        fc1_weights[59][22] = 16'sd-9;
        fc1_weights[59][23] = 16'sd-2;
        fc1_weights[59][24] = 16'sd1;
        fc1_weights[59][25] = 16'sd-29;
        fc1_weights[59][26] = 16'sd-51;
        fc1_weights[59][27] = 16'sd-40;
        fc1_weights[59][28] = 16'sd-49;
        fc1_weights[59][29] = 16'sd-18;
        fc1_weights[59][30] = 16'sd6;
        fc1_weights[59][31] = 16'sd24;
        fc1_weights[59][32] = 16'sd23;
        fc1_weights[59][33] = 16'sd47;
        fc1_weights[59][34] = 16'sd3;
        fc1_weights[59][35] = 16'sd-2;
        fc1_weights[59][36] = 16'sd53;
        fc1_weights[59][37] = 16'sd54;
        fc1_weights[59][38] = 16'sd8;
        fc1_weights[59][39] = 16'sd-69;
        fc1_weights[59][40] = 16'sd51;
        fc1_weights[59][41] = 16'sd27;
        fc1_weights[59][42] = 16'sd-38;
        fc1_weights[59][43] = 16'sd5;
        fc1_weights[59][44] = 16'sd25;
        fc1_weights[59][45] = 16'sd-42;
        fc1_weights[59][46] = 16'sd-21;
        fc1_weights[59][47] = 16'sd3;
        fc1_weights[59][48] = 16'sd39;
        fc1_weights[59][49] = 16'sd8;
        fc1_weights[59][50] = 16'sd-42;
        fc1_weights[59][51] = 16'sd-43;
        fc1_weights[59][52] = 16'sd-32;
        fc1_weights[59][53] = 16'sd-27;
        fc1_weights[59][54] = 16'sd-32;
        fc1_weights[59][55] = 16'sd-18;
        fc1_weights[59][56] = 16'sd-9;
        fc1_weights[59][57] = 16'sd10;
        fc1_weights[59][58] = 16'sd4;
        fc1_weights[59][59] = 16'sd8;
        fc1_weights[59][60] = 16'sd16;
        fc1_weights[59][61] = 16'sd2;
        fc1_weights[59][62] = 16'sd-9;
        fc1_weights[59][63] = 16'sd-13;
        fc1_weights[59][64] = 16'sd-5;
        fc1_weights[59][65] = 16'sd-19;
        fc1_weights[59][66] = 16'sd9;
        fc1_weights[59][67] = 16'sd-40;
        fc1_weights[59][68] = 16'sd-22;
        fc1_weights[59][69] = 16'sd-7;
        fc1_weights[59][70] = 16'sd-51;
        fc1_weights[59][71] = 16'sd-5;
        fc1_weights[59][72] = 16'sd12;
        fc1_weights[59][73] = 16'sd-12;
        fc1_weights[59][74] = 16'sd-30;
        fc1_weights[59][75] = 16'sd-51;
        fc1_weights[59][76] = 16'sd-35;
        fc1_weights[59][77] = 16'sd-64;
        fc1_weights[59][78] = 16'sd-26;
        fc1_weights[59][79] = 16'sd-3;
        fc1_weights[59][80] = 16'sd-41;
        fc1_weights[59][81] = 16'sd16;
        fc1_weights[59][82] = 16'sd13;
        fc1_weights[59][83] = 16'sd26;
        fc1_weights[59][84] = 16'sd-3;
        fc1_weights[59][85] = 16'sd-34;
        fc1_weights[59][86] = 16'sd-42;
        fc1_weights[59][87] = 16'sd-56;
        fc1_weights[59][88] = 16'sd-70;
        fc1_weights[59][89] = 16'sd135;
        fc1_weights[59][90] = 16'sd8;
        fc1_weights[59][91] = 16'sd64;
        fc1_weights[59][92] = 16'sd32;
        fc1_weights[59][93] = 16'sd62;
        fc1_weights[59][94] = 16'sd20;
        fc1_weights[59][95] = 16'sd25;
        fc1_weights[59][96] = 16'sd-21;
        fc1_weights[59][97] = 16'sd-54;
        fc1_weights[59][98] = 16'sd-33;
        fc1_weights[59][99] = 16'sd-37;
        fc1_weights[59][100] = 16'sd-4;
        fc1_weights[59][101] = 16'sd-44;
        fc1_weights[59][102] = 16'sd-27;
        fc1_weights[59][103] = 16'sd-46;
        fc1_weights[59][104] = 16'sd-28;
        fc1_weights[59][105] = 16'sd-25;
        fc1_weights[59][106] = 16'sd-47;
        fc1_weights[59][107] = 16'sd-36;
        fc1_weights[59][108] = 16'sd-16;
        fc1_weights[59][109] = 16'sd35;
        fc1_weights[59][110] = 16'sd9;
        fc1_weights[59][111] = 16'sd-29;
        fc1_weights[59][112] = 16'sd18;
        fc1_weights[59][113] = 16'sd19;
        fc1_weights[59][114] = 16'sd39;
        fc1_weights[59][115] = 16'sd-1;
        fc1_weights[59][116] = 16'sd27;
        fc1_weights[59][117] = 16'sd59;
        fc1_weights[59][118] = 16'sd-16;
        fc1_weights[59][119] = 16'sd45;
        fc1_weights[59][120] = 16'sd31;
        fc1_weights[59][121] = 16'sd-10;
        fc1_weights[59][122] = 16'sd34;
        fc1_weights[59][123] = 16'sd-8;
        fc1_weights[59][124] = 16'sd2;
        fc1_weights[59][125] = 16'sd-43;
        fc1_weights[59][126] = 16'sd-53;
        fc1_weights[59][127] = 16'sd-55;
        fc1_weights[59][128] = 16'sd-51;
        fc1_weights[59][129] = 16'sd-83;
        fc1_weights[59][130] = 16'sd-23;
        fc1_weights[59][131] = 16'sd-41;
        fc1_weights[59][132] = 16'sd-21;
        fc1_weights[59][133] = 16'sd1;
        fc1_weights[59][134] = 16'sd8;
        fc1_weights[59][135] = 16'sd48;
        fc1_weights[59][136] = 16'sd6;
        fc1_weights[59][137] = 16'sd28;
        fc1_weights[59][138] = 16'sd-15;
        fc1_weights[59][139] = 16'sd69;
        fc1_weights[59][140] = 16'sd68;
        fc1_weights[59][141] = 16'sd-23;
        fc1_weights[59][142] = 16'sd43;
        fc1_weights[59][143] = 16'sd53;
        fc1_weights[59][144] = 16'sd46;
        fc1_weights[59][145] = 16'sd1;
        fc1_weights[59][146] = 16'sd7;
        fc1_weights[59][147] = 16'sd45;
        fc1_weights[59][148] = 16'sd60;
        fc1_weights[59][149] = 16'sd23;
        fc1_weights[59][150] = 16'sd-30;
        fc1_weights[59][151] = 16'sd-15;
        fc1_weights[59][152] = 16'sd9;
        fc1_weights[59][153] = 16'sd-10;
        fc1_weights[59][154] = 16'sd-10;
        fc1_weights[59][155] = 16'sd43;
        fc1_weights[59][156] = 16'sd2;
        fc1_weights[59][157] = 16'sd-30;
        fc1_weights[59][158] = 16'sd-18;
        fc1_weights[59][159] = 16'sd24;
        fc1_weights[59][160] = 16'sd-34;
        fc1_weights[59][161] = 16'sd-76;
        fc1_weights[59][162] = 16'sd-20;
        fc1_weights[59][163] = 16'sd-8;
        fc1_weights[59][164] = 16'sd14;
        fc1_weights[59][165] = 16'sd18;
        fc1_weights[59][166] = 16'sd48;
        fc1_weights[59][167] = 16'sd16;
        fc1_weights[59][168] = 16'sd15;
        fc1_weights[59][169] = 16'sd-48;
        fc1_weights[59][170] = 16'sd-3;
        fc1_weights[59][171] = 16'sd18;
        fc1_weights[59][172] = 16'sd22;
        fc1_weights[59][173] = 16'sd21;
        fc1_weights[59][174] = 16'sd35;
        fc1_weights[59][175] = 16'sd103;
        fc1_weights[59][176] = 16'sd53;
        fc1_weights[59][177] = 16'sd-4;
        fc1_weights[59][178] = 16'sd11;
        fc1_weights[59][179] = 16'sd40;
        fc1_weights[59][180] = 16'sd20;
        fc1_weights[59][181] = 16'sd7;
        fc1_weights[59][182] = 16'sd-19;
        fc1_weights[59][183] = 16'sd28;
        fc1_weights[59][184] = 16'sd-18;
        fc1_weights[59][185] = 16'sd55;
        fc1_weights[59][186] = 16'sd-48;
        fc1_weights[59][187] = 16'sd-12;
        fc1_weights[59][188] = 16'sd-3;
        fc1_weights[59][189] = 16'sd17;
        fc1_weights[59][190] = 16'sd44;
        fc1_weights[59][191] = 16'sd16;
        fc1_weights[59][192] = 16'sd-13;
        fc1_weights[59][193] = 16'sd12;
        fc1_weights[59][194] = 16'sd0;
        fc1_weights[59][195] = 16'sd-30;
        fc1_weights[59][196] = 16'sd-30;
        fc1_weights[59][197] = 16'sd32;
        fc1_weights[59][198] = 16'sd-22;
        fc1_weights[59][199] = 16'sd11;
        fc1_weights[59][200] = 16'sd-30;
        fc1_weights[59][201] = 16'sd22;
        fc1_weights[59][202] = 16'sd-4;
        fc1_weights[59][203] = 16'sd23;
        fc1_weights[59][204] = 16'sd42;
        fc1_weights[59][205] = 16'sd64;
        fc1_weights[59][206] = 16'sd-33;
        fc1_weights[59][207] = 16'sd-9;
        fc1_weights[60][0] = 16'sd-35;
        fc1_weights[60][1] = 16'sd39;
        fc1_weights[60][2] = 16'sd-13;
        fc1_weights[60][3] = 16'sd-23;
        fc1_weights[60][4] = 16'sd-50;
        fc1_weights[60][5] = 16'sd-18;
        fc1_weights[60][6] = 16'sd-6;
        fc1_weights[60][7] = 16'sd36;
        fc1_weights[60][8] = 16'sd-16;
        fc1_weights[60][9] = 16'sd-8;
        fc1_weights[60][10] = 16'sd42;
        fc1_weights[60][11] = 16'sd97;
        fc1_weights[60][12] = 16'sd-1;
        fc1_weights[60][13] = 16'sd-30;
        fc1_weights[60][14] = 16'sd-75;
        fc1_weights[60][15] = 16'sd-20;
        fc1_weights[60][16] = 16'sd-23;
        fc1_weights[60][17] = 16'sd-32;
        fc1_weights[60][18] = 16'sd-18;
        fc1_weights[60][19] = 16'sd-57;
        fc1_weights[60][20] = 16'sd5;
        fc1_weights[60][21] = 16'sd55;
        fc1_weights[60][22] = 16'sd-44;
        fc1_weights[60][23] = 16'sd-34;
        fc1_weights[60][24] = 16'sd6;
        fc1_weights[60][25] = 16'sd27;
        fc1_weights[60][26] = 16'sd-51;
        fc1_weights[60][27] = 16'sd-16;
        fc1_weights[60][28] = 16'sd-9;
        fc1_weights[60][29] = 16'sd15;
        fc1_weights[60][30] = 16'sd-26;
        fc1_weights[60][31] = 16'sd-17;
        fc1_weights[60][32] = 16'sd-17;
        fc1_weights[60][33] = 16'sd-44;
        fc1_weights[60][34] = 16'sd3;
        fc1_weights[60][35] = 16'sd11;
        fc1_weights[60][36] = 16'sd32;
        fc1_weights[60][37] = 16'sd67;
        fc1_weights[60][38] = 16'sd84;
        fc1_weights[60][39] = 16'sd5;
        fc1_weights[60][40] = 16'sd18;
        fc1_weights[60][41] = 16'sd-96;
        fc1_weights[60][42] = 16'sd-50;
        fc1_weights[60][43] = 16'sd7;
        fc1_weights[60][44] = 16'sd24;
        fc1_weights[60][45] = 16'sd17;
        fc1_weights[60][46] = 16'sd59;
        fc1_weights[60][47] = 16'sd1;
        fc1_weights[60][48] = 16'sd33;
        fc1_weights[60][49] = 16'sd47;
        fc1_weights[60][50] = 16'sd-30;
        fc1_weights[60][51] = 16'sd-41;
        fc1_weights[60][52] = 16'sd-61;
        fc1_weights[60][53] = 16'sd-42;
        fc1_weights[60][54] = 16'sd-14;
        fc1_weights[60][55] = 16'sd3;
        fc1_weights[60][56] = 16'sd40;
        fc1_weights[60][57] = 16'sd5;
        fc1_weights[60][58] = 16'sd-45;
        fc1_weights[60][59] = 16'sd-57;
        fc1_weights[60][60] = 16'sd50;
        fc1_weights[60][61] = 16'sd4;
        fc1_weights[60][62] = 16'sd4;
        fc1_weights[60][63] = 16'sd73;
        fc1_weights[60][64] = 16'sd137;
        fc1_weights[60][65] = 16'sd-66;
        fc1_weights[60][66] = 16'sd-92;
        fc1_weights[60][67] = 16'sd-27;
        fc1_weights[60][68] = 16'sd-39;
        fc1_weights[60][69] = 16'sd60;
        fc1_weights[60][70] = 16'sd64;
        fc1_weights[60][71] = 16'sd15;
        fc1_weights[60][72] = 16'sd38;
        fc1_weights[60][73] = 16'sd43;
        fc1_weights[60][74] = 16'sd88;
        fc1_weights[60][75] = 16'sd-20;
        fc1_weights[60][76] = 16'sd6;
        fc1_weights[60][77] = 16'sd29;
        fc1_weights[60][78] = 16'sd-25;
        fc1_weights[60][79] = 16'sd7;
        fc1_weights[60][80] = 16'sd-12;
        fc1_weights[60][81] = 16'sd15;
        fc1_weights[60][82] = 16'sd-13;
        fc1_weights[60][83] = 16'sd-33;
        fc1_weights[60][84] = 16'sd27;
        fc1_weights[60][85] = 16'sd-59;
        fc1_weights[60][86] = 16'sd-8;
        fc1_weights[60][87] = 16'sd55;
        fc1_weights[60][88] = 16'sd46;
        fc1_weights[60][89] = 16'sd-58;
        fc1_weights[60][90] = 16'sd102;
        fc1_weights[60][91] = 16'sd26;
        fc1_weights[60][92] = 16'sd49;
        fc1_weights[60][93] = 16'sd-44;
        fc1_weights[60][94] = 16'sd-18;
        fc1_weights[60][95] = 16'sd28;
        fc1_weights[60][96] = 16'sd5;
        fc1_weights[60][97] = 16'sd-8;
        fc1_weights[60][98] = 16'sd-1;
        fc1_weights[60][99] = 16'sd-15;
        fc1_weights[60][100] = 16'sd13;
        fc1_weights[60][101] = 16'sd68;
        fc1_weights[60][102] = 16'sd-49;
        fc1_weights[60][103] = 16'sd15;
        fc1_weights[60][104] = 16'sd5;
        fc1_weights[60][105] = 16'sd-111;
        fc1_weights[60][106] = 16'sd-14;
        fc1_weights[60][107] = 16'sd9;
        fc1_weights[60][108] = 16'sd-55;
        fc1_weights[60][109] = 16'sd-50;
        fc1_weights[60][110] = 16'sd8;
        fc1_weights[60][111] = 16'sd-25;
        fc1_weights[60][112] = 16'sd85;
        fc1_weights[60][113] = 16'sd2;
        fc1_weights[60][114] = 16'sd-52;
        fc1_weights[60][115] = 16'sd-13;
        fc1_weights[60][116] = 16'sd46;
        fc1_weights[60][117] = 16'sd-31;
        fc1_weights[60][118] = 16'sd46;
        fc1_weights[60][119] = 16'sd7;
        fc1_weights[60][120] = 16'sd-20;
        fc1_weights[60][121] = 16'sd21;
        fc1_weights[60][122] = 16'sd-18;
        fc1_weights[60][123] = 16'sd-13;
        fc1_weights[60][124] = 16'sd-1;
        fc1_weights[60][125] = 16'sd41;
        fc1_weights[60][126] = 16'sd56;
        fc1_weights[60][127] = 16'sd61;
        fc1_weights[60][128] = 16'sd2;
        fc1_weights[60][129] = 16'sd-5;
        fc1_weights[60][130] = 16'sd-31;
        fc1_weights[60][131] = 16'sd-5;
        fc1_weights[60][132] = 16'sd28;
        fc1_weights[60][133] = 16'sd-10;
        fc1_weights[60][134] = 16'sd-4;
        fc1_weights[60][135] = 16'sd9;
        fc1_weights[60][136] = 16'sd36;
        fc1_weights[60][137] = 16'sd-24;
        fc1_weights[60][138] = 16'sd138;
        fc1_weights[60][139] = 16'sd33;
        fc1_weights[60][140] = 16'sd-44;
        fc1_weights[60][141] = 16'sd-11;
        fc1_weights[60][142] = 16'sd-25;
        fc1_weights[60][143] = 16'sd-53;
        fc1_weights[60][144] = 16'sd11;
        fc1_weights[60][145] = 16'sd31;
        fc1_weights[60][146] = 16'sd68;
        fc1_weights[60][147] = 16'sd-35;
        fc1_weights[60][148] = 16'sd-23;
        fc1_weights[60][149] = 16'sd44;
        fc1_weights[60][150] = 16'sd44;
        fc1_weights[60][151] = 16'sd93;
        fc1_weights[60][152] = 16'sd18;
        fc1_weights[60][153] = 16'sd-1;
        fc1_weights[60][154] = 16'sd-22;
        fc1_weights[60][155] = 16'sd5;
        fc1_weights[60][156] = 16'sd-12;
        fc1_weights[60][157] = 16'sd-58;
        fc1_weights[60][158] = 16'sd-12;
        fc1_weights[60][159] = 16'sd40;
        fc1_weights[60][160] = 16'sd-35;
        fc1_weights[60][161] = 16'sd-28;
        fc1_weights[60][162] = 16'sd108;
        fc1_weights[60][163] = 16'sd18;
        fc1_weights[60][164] = 16'sd20;
        fc1_weights[60][165] = 16'sd-81;
        fc1_weights[60][166] = 16'sd9;
        fc1_weights[60][167] = 16'sd-1;
        fc1_weights[60][168] = 16'sd9;
        fc1_weights[60][169] = 16'sd-57;
        fc1_weights[60][170] = 16'sd24;
        fc1_weights[60][171] = 16'sd-99;
        fc1_weights[60][172] = 16'sd-12;
        fc1_weights[60][173] = 16'sd-5;
        fc1_weights[60][174] = 16'sd-18;
        fc1_weights[60][175] = 16'sd-45;
        fc1_weights[60][176] = 16'sd-37;
        fc1_weights[60][177] = 16'sd45;
        fc1_weights[60][178] = 16'sd-5;
        fc1_weights[60][179] = 16'sd40;
        fc1_weights[60][180] = 16'sd8;
        fc1_weights[60][181] = 16'sd63;
        fc1_weights[60][182] = 16'sd60;
        fc1_weights[60][183] = 16'sd-3;
        fc1_weights[60][184] = 16'sd15;
        fc1_weights[60][185] = 16'sd87;
        fc1_weights[60][186] = 16'sd23;
        fc1_weights[60][187] = 16'sd11;
        fc1_weights[60][188] = 16'sd40;
        fc1_weights[60][189] = 16'sd-8;
        fc1_weights[60][190] = 16'sd-5;
        fc1_weights[60][191] = 16'sd13;
        fc1_weights[60][192] = 16'sd-55;
        fc1_weights[60][193] = 16'sd-31;
        fc1_weights[60][194] = 16'sd-38;
        fc1_weights[60][195] = 16'sd-2;
        fc1_weights[60][196] = 16'sd-43;
        fc1_weights[60][197] = 16'sd78;
        fc1_weights[60][198] = 16'sd-45;
        fc1_weights[60][199] = 16'sd-47;
        fc1_weights[60][200] = 16'sd15;
        fc1_weights[60][201] = 16'sd-3;
        fc1_weights[60][202] = 16'sd-52;
        fc1_weights[60][203] = 16'sd17;
        fc1_weights[60][204] = 16'sd11;
        fc1_weights[60][205] = 16'sd4;
        fc1_weights[60][206] = 16'sd-28;
        fc1_weights[60][207] = 16'sd68;
        fc1_weights[61][0] = 16'sd-23;
        fc1_weights[61][1] = 16'sd2;
        fc1_weights[61][2] = 16'sd36;
        fc1_weights[61][3] = 16'sd77;
        fc1_weights[61][4] = 16'sd42;
        fc1_weights[61][5] = 16'sd55;
        fc1_weights[61][6] = 16'sd50;
        fc1_weights[61][7] = 16'sd78;
        fc1_weights[61][8] = 16'sd58;
        fc1_weights[61][9] = 16'sd33;
        fc1_weights[61][10] = 16'sd41;
        fc1_weights[61][11] = 16'sd11;
        fc1_weights[61][12] = 16'sd20;
        fc1_weights[61][13] = 16'sd8;
        fc1_weights[61][14] = 16'sd-9;
        fc1_weights[61][15] = 16'sd-21;
        fc1_weights[61][16] = 16'sd-17;
        fc1_weights[61][17] = 16'sd-41;
        fc1_weights[61][18] = 16'sd-11;
        fc1_weights[61][19] = 16'sd-25;
        fc1_weights[61][20] = 16'sd19;
        fc1_weights[61][21] = 16'sd19;
        fc1_weights[61][22] = 16'sd29;
        fc1_weights[61][23] = 16'sd28;
        fc1_weights[61][24] = 16'sd46;
        fc1_weights[61][25] = 16'sd49;
        fc1_weights[61][26] = 16'sd-21;
        fc1_weights[61][27] = 16'sd6;
        fc1_weights[61][28] = 16'sd10;
        fc1_weights[61][29] = 16'sd67;
        fc1_weights[61][30] = 16'sd39;
        fc1_weights[61][31] = 16'sd26;
        fc1_weights[61][32] = 16'sd45;
        fc1_weights[61][33] = 16'sd69;
        fc1_weights[61][34] = 16'sd60;
        fc1_weights[61][35] = 16'sd35;
        fc1_weights[61][36] = 16'sd37;
        fc1_weights[61][37] = 16'sd53;
        fc1_weights[61][38] = 16'sd34;
        fc1_weights[61][39] = 16'sd1;
        fc1_weights[61][40] = 16'sd9;
        fc1_weights[61][41] = 16'sd-11;
        fc1_weights[61][42] = 16'sd-6;
        fc1_weights[61][43] = 16'sd-3;
        fc1_weights[61][44] = 16'sd-5;
        fc1_weights[61][45] = 16'sd26;
        fc1_weights[61][46] = 16'sd15;
        fc1_weights[61][47] = 16'sd52;
        fc1_weights[61][48] = 16'sd37;
        fc1_weights[61][49] = 16'sd69;
        fc1_weights[61][50] = 16'sd22;
        fc1_weights[61][51] = 16'sd38;
        fc1_weights[61][52] = 16'sd-12;
        fc1_weights[61][53] = 16'sd-31;
        fc1_weights[61][54] = 16'sd14;
        fc1_weights[61][55] = 16'sd29;
        fc1_weights[61][56] = 16'sd54;
        fc1_weights[61][57] = 16'sd-27;
        fc1_weights[61][58] = 16'sd-9;
        fc1_weights[61][59] = 16'sd18;
        fc1_weights[61][60] = 16'sd0;
        fc1_weights[61][61] = 16'sd-33;
        fc1_weights[61][62] = 16'sd30;
        fc1_weights[61][63] = 16'sd18;
        fc1_weights[61][64] = 16'sd-1;
        fc1_weights[61][65] = 16'sd15;
        fc1_weights[61][66] = 16'sd-17;
        fc1_weights[61][67] = 16'sd3;
        fc1_weights[61][68] = 16'sd6;
        fc1_weights[61][69] = 16'sd64;
        fc1_weights[61][70] = 16'sd29;
        fc1_weights[61][71] = 16'sd65;
        fc1_weights[61][72] = 16'sd71;
        fc1_weights[61][73] = 16'sd81;
        fc1_weights[61][74] = 16'sd70;
        fc1_weights[61][75] = 16'sd61;
        fc1_weights[61][76] = 16'sd3;
        fc1_weights[61][77] = 16'sd24;
        fc1_weights[61][78] = 16'sd-30;
        fc1_weights[61][79] = 16'sd-3;
        fc1_weights[61][80] = 16'sd30;
        fc1_weights[61][81] = 16'sd20;
        fc1_weights[61][82] = 16'sd7;
        fc1_weights[61][83] = 16'sd31;
        fc1_weights[61][84] = 16'sd25;
        fc1_weights[61][85] = 16'sd37;
        fc1_weights[61][86] = 16'sd22;
        fc1_weights[61][87] = 16'sd26;
        fc1_weights[61][88] = 16'sd5;
        fc1_weights[61][89] = 16'sd36;
        fc1_weights[61][90] = 16'sd-71;
        fc1_weights[61][91] = 16'sd-50;
        fc1_weights[61][92] = 16'sd-36;
        fc1_weights[61][93] = 16'sd2;
        fc1_weights[61][94] = 16'sd-18;
        fc1_weights[61][95] = 16'sd-5;
        fc1_weights[61][96] = 16'sd9;
        fc1_weights[61][97] = 16'sd0;
        fc1_weights[61][98] = 16'sd20;
        fc1_weights[61][99] = 16'sd25;
        fc1_weights[61][100] = 16'sd40;
        fc1_weights[61][101] = 16'sd49;
        fc1_weights[61][102] = 16'sd1;
        fc1_weights[61][103] = 16'sd-22;
        fc1_weights[61][104] = 16'sd-44;
        fc1_weights[61][105] = 16'sd-31;
        fc1_weights[61][106] = 16'sd-11;
        fc1_weights[61][107] = 16'sd5;
        fc1_weights[61][108] = 16'sd12;
        fc1_weights[61][109] = 16'sd25;
        fc1_weights[61][110] = 16'sd-6;
        fc1_weights[61][111] = 16'sd0;
        fc1_weights[61][112] = 16'sd-9;
        fc1_weights[61][113] = 16'sd18;
        fc1_weights[61][114] = 16'sd-41;
        fc1_weights[61][115] = 16'sd-33;
        fc1_weights[61][116] = 16'sd3;
        fc1_weights[61][117] = 16'sd7;
        fc1_weights[61][118] = 16'sd16;
        fc1_weights[61][119] = 16'sd-11;
        fc1_weights[61][120] = 16'sd-42;
        fc1_weights[61][121] = 16'sd-14;
        fc1_weights[61][122] = 16'sd18;
        fc1_weights[61][123] = 16'sd-10;
        fc1_weights[61][124] = 16'sd26;
        fc1_weights[61][125] = 16'sd33;
        fc1_weights[61][126] = 16'sd36;
        fc1_weights[61][127] = 16'sd-11;
        fc1_weights[61][128] = 16'sd0;
        fc1_weights[61][129] = 16'sd4;
        fc1_weights[61][130] = 16'sd1;
        fc1_weights[61][131] = 16'sd44;
        fc1_weights[61][132] = 16'sd19;
        fc1_weights[61][133] = 16'sd-33;
        fc1_weights[61][134] = 16'sd15;
        fc1_weights[61][135] = 16'sd22;
        fc1_weights[61][136] = 16'sd25;
        fc1_weights[61][137] = 16'sd36;
        fc1_weights[61][138] = 16'sd-22;
        fc1_weights[61][139] = 16'sd23;
        fc1_weights[61][140] = 16'sd-32;
        fc1_weights[61][141] = 16'sd-28;
        fc1_weights[61][142] = 16'sd7;
        fc1_weights[61][143] = 16'sd35;
        fc1_weights[61][144] = 16'sd8;
        fc1_weights[61][145] = 16'sd22;
        fc1_weights[61][146] = 16'sd-19;
        fc1_weights[61][147] = 16'sd-28;
        fc1_weights[61][148] = 16'sd-24;
        fc1_weights[61][149] = 16'sd-46;
        fc1_weights[61][150] = 16'sd2;
        fc1_weights[61][151] = 16'sd-9;
        fc1_weights[61][152] = 16'sd-6;
        fc1_weights[61][153] = 16'sd-16;
        fc1_weights[61][154] = 16'sd-47;
        fc1_weights[61][155] = 16'sd-26;
        fc1_weights[61][156] = 16'sd-9;
        fc1_weights[61][157] = 16'sd-13;
        fc1_weights[61][158] = 16'sd27;
        fc1_weights[61][159] = 16'sd40;
        fc1_weights[61][160] = 16'sd37;
        fc1_weights[61][161] = 16'sd3;
        fc1_weights[61][162] = 16'sd-24;
        fc1_weights[61][163] = 16'sd-5;
        fc1_weights[61][164] = 16'sd13;
        fc1_weights[61][165] = 16'sd2;
        fc1_weights[61][166] = 16'sd20;
        fc1_weights[61][167] = 16'sd8;
        fc1_weights[61][168] = 16'sd10;
        fc1_weights[61][169] = 16'sd9;
        fc1_weights[61][170] = 16'sd-21;
        fc1_weights[61][171] = 16'sd5;
        fc1_weights[61][172] = 16'sd9;
        fc1_weights[61][173] = 16'sd-21;
        fc1_weights[61][174] = 16'sd2;
        fc1_weights[61][175] = 16'sd-19;
        fc1_weights[61][176] = 16'sd-10;
        fc1_weights[61][177] = 16'sd-17;
        fc1_weights[61][178] = 16'sd7;
        fc1_weights[61][179] = 16'sd-18;
        fc1_weights[61][180] = 16'sd-27;
        fc1_weights[61][181] = 16'sd1;
        fc1_weights[61][182] = 16'sd1;
        fc1_weights[61][183] = 16'sd25;
        fc1_weights[61][184] = 16'sd22;
        fc1_weights[61][185] = 16'sd9;
        fc1_weights[61][186] = 16'sd-3;
        fc1_weights[61][187] = 16'sd10;
        fc1_weights[61][188] = 16'sd27;
        fc1_weights[61][189] = 16'sd16;
        fc1_weights[61][190] = 16'sd-6;
        fc1_weights[61][191] = 16'sd-2;
        fc1_weights[61][192] = 16'sd22;
        fc1_weights[61][193] = 16'sd23;
        fc1_weights[61][194] = 16'sd8;
        fc1_weights[61][195] = 16'sd-9;
        fc1_weights[61][196] = 16'sd-16;
        fc1_weights[61][197] = 16'sd-14;
        fc1_weights[61][198] = 16'sd26;
        fc1_weights[61][199] = 16'sd-39;
        fc1_weights[61][200] = 16'sd-1;
        fc1_weights[61][201] = 16'sd-4;
        fc1_weights[61][202] = 16'sd19;
        fc1_weights[61][203] = 16'sd-6;
        fc1_weights[61][204] = 16'sd-16;
        fc1_weights[61][205] = 16'sd-30;
        fc1_weights[61][206] = 16'sd2;
        fc1_weights[61][207] = 16'sd-11;
        fc1_weights[62][0] = 16'sd41;
        fc1_weights[62][1] = 16'sd-13;
        fc1_weights[62][2] = 16'sd-42;
        fc1_weights[62][3] = 16'sd-49;
        fc1_weights[62][4] = 16'sd5;
        fc1_weights[62][5] = 16'sd55;
        fc1_weights[62][6] = 16'sd18;
        fc1_weights[62][7] = 16'sd-1;
        fc1_weights[62][8] = 16'sd-28;
        fc1_weights[62][9] = 16'sd-24;
        fc1_weights[62][10] = 16'sd-41;
        fc1_weights[62][11] = 16'sd-50;
        fc1_weights[62][12] = 16'sd-37;
        fc1_weights[62][13] = 16'sd16;
        fc1_weights[62][14] = 16'sd-18;
        fc1_weights[62][15] = 16'sd27;
        fc1_weights[62][16] = 16'sd-5;
        fc1_weights[62][17] = 16'sd-84;
        fc1_weights[62][18] = 16'sd-45;
        fc1_weights[62][19] = 16'sd-20;
        fc1_weights[62][20] = 16'sd16;
        fc1_weights[62][21] = 16'sd-98;
        fc1_weights[62][22] = 16'sd-29;
        fc1_weights[62][23] = 16'sd-18;
        fc1_weights[62][24] = 16'sd23;
        fc1_weights[62][25] = 16'sd-52;
        fc1_weights[62][26] = 16'sd-37;
        fc1_weights[62][27] = 16'sd-25;
        fc1_weights[62][28] = 16'sd-9;
        fc1_weights[62][29] = 16'sd2;
        fc1_weights[62][30] = 16'sd-32;
        fc1_weights[62][31] = 16'sd55;
        fc1_weights[62][32] = 16'sd19;
        fc1_weights[62][33] = 16'sd3;
        fc1_weights[62][34] = 16'sd-39;
        fc1_weights[62][35] = 16'sd-11;
        fc1_weights[62][36] = 16'sd-2;
        fc1_weights[62][37] = 16'sd-74;
        fc1_weights[62][38] = 16'sd-29;
        fc1_weights[62][39] = 16'sd6;
        fc1_weights[62][40] = 16'sd-2;
        fc1_weights[62][41] = 16'sd0;
        fc1_weights[62][42] = 16'sd-36;
        fc1_weights[62][43] = 16'sd-45;
        fc1_weights[62][44] = 16'sd-25;
        fc1_weights[62][45] = 16'sd-13;
        fc1_weights[62][46] = 16'sd4;
        fc1_weights[62][47] = 16'sd-48;
        fc1_weights[62][48] = 16'sd-24;
        fc1_weights[62][49] = 16'sd-38;
        fc1_weights[62][50] = 16'sd-37;
        fc1_weights[62][51] = 16'sd-10;
        fc1_weights[62][52] = 16'sd23;
        fc1_weights[62][53] = 16'sd-22;
        fc1_weights[62][54] = 16'sd-24;
        fc1_weights[62][55] = 16'sd-29;
        fc1_weights[62][56] = 16'sd5;
        fc1_weights[62][57] = 16'sd66;
        fc1_weights[62][58] = 16'sd14;
        fc1_weights[62][59] = 16'sd49;
        fc1_weights[62][60] = 16'sd96;
        fc1_weights[62][61] = 16'sd9;
        fc1_weights[62][62] = 16'sd-62;
        fc1_weights[62][63] = 16'sd-21;
        fc1_weights[62][64] = 16'sd-3;
        fc1_weights[62][65] = 16'sd21;
        fc1_weights[62][66] = 16'sd1;
        fc1_weights[62][67] = 16'sd-5;
        fc1_weights[62][68] = 16'sd-23;
        fc1_weights[62][69] = 16'sd-93;
        fc1_weights[62][70] = 16'sd14;
        fc1_weights[62][71] = 16'sd86;
        fc1_weights[62][72] = 16'sd76;
        fc1_weights[62][73] = 16'sd12;
        fc1_weights[62][74] = 16'sd27;
        fc1_weights[62][75] = 16'sd-34;
        fc1_weights[62][76] = 16'sd36;
        fc1_weights[62][77] = 16'sd-20;
        fc1_weights[62][78] = 16'sd6;
        fc1_weights[62][79] = 16'sd34;
        fc1_weights[62][80] = 16'sd-33;
        fc1_weights[62][81] = 16'sd4;
        fc1_weights[62][82] = 16'sd-6;
        fc1_weights[62][83] = 16'sd48;
        fc1_weights[62][84] = 16'sd-54;
        fc1_weights[62][85] = 16'sd31;
        fc1_weights[62][86] = 16'sd83;
        fc1_weights[62][87] = 16'sd34;
        fc1_weights[62][88] = 16'sd39;
        fc1_weights[62][89] = 16'sd-14;
        fc1_weights[62][90] = 16'sd54;
        fc1_weights[62][91] = 16'sd10;
        fc1_weights[62][92] = 16'sd-53;
        fc1_weights[62][93] = 16'sd-63;
        fc1_weights[62][94] = 16'sd-108;
        fc1_weights[62][95] = 16'sd-23;
        fc1_weights[62][96] = 16'sd-4;
        fc1_weights[62][97] = 16'sd19;
        fc1_weights[62][98] = 16'sd14;
        fc1_weights[62][99] = 16'sd-16;
        fc1_weights[62][100] = 16'sd16;
        fc1_weights[62][101] = 16'sd-93;
        fc1_weights[62][102] = 16'sd-35;
        fc1_weights[62][103] = 16'sd-12;
        fc1_weights[62][104] = 16'sd43;
        fc1_weights[62][105] = 16'sd-39;
        fc1_weights[62][106] = 16'sd6;
        fc1_weights[62][107] = 16'sd40;
        fc1_weights[62][108] = 16'sd18;
        fc1_weights[62][109] = 16'sd52;
        fc1_weights[62][110] = 16'sd24;
        fc1_weights[62][111] = 16'sd8;
        fc1_weights[62][112] = 16'sd112;
        fc1_weights[62][113] = 16'sd69;
        fc1_weights[62][114] = 16'sd9;
        fc1_weights[62][115] = 16'sd-26;
        fc1_weights[62][116] = 16'sd8;
        fc1_weights[62][117] = 16'sd-16;
        fc1_weights[62][118] = 16'sd5;
        fc1_weights[62][119] = 16'sd47;
        fc1_weights[62][120] = 16'sd-14;
        fc1_weights[62][121] = 16'sd-4;
        fc1_weights[62][122] = 16'sd-12;
        fc1_weights[62][123] = 16'sd-17;
        fc1_weights[62][124] = 16'sd-14;
        fc1_weights[62][125] = 16'sd11;
        fc1_weights[62][126] = 16'sd-38;
        fc1_weights[62][127] = 16'sd-23;
        fc1_weights[62][128] = 16'sd3;
        fc1_weights[62][129] = 16'sd-38;
        fc1_weights[62][130] = 16'sd67;
        fc1_weights[62][131] = 16'sd93;
        fc1_weights[62][132] = 16'sd68;
        fc1_weights[62][133] = 16'sd40;
        fc1_weights[62][134] = 16'sd-10;
        fc1_weights[62][135] = 16'sd32;
        fc1_weights[62][136] = 16'sd18;
        fc1_weights[62][137] = 16'sd-6;
        fc1_weights[62][138] = 16'sd9;
        fc1_weights[62][139] = 16'sd13;
        fc1_weights[62][140] = 16'sd-1;
        fc1_weights[62][141] = 16'sd-75;
        fc1_weights[62][142] = 16'sd17;
        fc1_weights[62][143] = 16'sd13;
        fc1_weights[62][144] = 16'sd-15;
        fc1_weights[62][145] = 16'sd-16;
        fc1_weights[62][146] = 16'sd-42;
        fc1_weights[62][147] = 16'sd-16;
        fc1_weights[62][148] = 16'sd-34;
        fc1_weights[62][149] = 16'sd-61;
        fc1_weights[62][150] = 16'sd-63;
        fc1_weights[62][151] = 16'sd40;
        fc1_weights[62][152] = 16'sd-26;
        fc1_weights[62][153] = 16'sd-18;
        fc1_weights[62][154] = 16'sd-24;
        fc1_weights[62][155] = 16'sd8;
        fc1_weights[62][156] = 16'sd39;
        fc1_weights[62][157] = 16'sd17;
        fc1_weights[62][158] = 16'sd-6;
        fc1_weights[62][159] = 16'sd-16;
        fc1_weights[62][160] = 16'sd-44;
        fc1_weights[62][161] = 16'sd12;
        fc1_weights[62][162] = 16'sd-31;
        fc1_weights[62][163] = 16'sd0;
        fc1_weights[62][164] = 16'sd-11;
        fc1_weights[62][165] = 16'sd-63;
        fc1_weights[62][166] = 16'sd8;
        fc1_weights[62][167] = 16'sd-11;
        fc1_weights[62][168] = 16'sd-51;
        fc1_weights[62][169] = 16'sd12;
        fc1_weights[62][170] = 16'sd35;
        fc1_weights[62][171] = 16'sd-12;
        fc1_weights[62][172] = 16'sd-56;
        fc1_weights[62][173] = 16'sd1;
        fc1_weights[62][174] = 16'sd-32;
        fc1_weights[62][175] = 16'sd25;
        fc1_weights[62][176] = 16'sd-10;
        fc1_weights[62][177] = 16'sd-39;
        fc1_weights[62][178] = 16'sd-9;
        fc1_weights[62][179] = 16'sd-8;
        fc1_weights[62][180] = 16'sd-2;
        fc1_weights[62][181] = 16'sd-5;
        fc1_weights[62][182] = 16'sd-35;
        fc1_weights[62][183] = 16'sd-1;
        fc1_weights[62][184] = 16'sd-13;
        fc1_weights[62][185] = 16'sd28;
        fc1_weights[62][186] = 16'sd-99;
        fc1_weights[62][187] = 16'sd-95;
        fc1_weights[62][188] = 16'sd-73;
        fc1_weights[62][189] = 16'sd24;
        fc1_weights[62][190] = 16'sd24;
        fc1_weights[62][191] = 16'sd0;
        fc1_weights[62][192] = 16'sd28;
        fc1_weights[62][193] = 16'sd4;
        fc1_weights[62][194] = 16'sd-1;
        fc1_weights[62][195] = 16'sd-6;
        fc1_weights[62][196] = 16'sd28;
        fc1_weights[62][197] = 16'sd71;
        fc1_weights[62][198] = 16'sd3;
        fc1_weights[62][199] = 16'sd5;
        fc1_weights[62][200] = 16'sd-1;
        fc1_weights[62][201] = 16'sd0;
        fc1_weights[62][202] = 16'sd-58;
        fc1_weights[62][203] = 16'sd-11;
        fc1_weights[62][204] = 16'sd-24;
        fc1_weights[62][205] = 16'sd-30;
        fc1_weights[62][206] = 16'sd-27;
        fc1_weights[62][207] = 16'sd8;
        fc1_weights[63][0] = 16'sd2;
        fc1_weights[63][1] = 16'sd4;
        fc1_weights[63][2] = 16'sd-29;
        fc1_weights[63][3] = 16'sd-17;
        fc1_weights[63][4] = 16'sd-38;
        fc1_weights[63][5] = 16'sd-15;
        fc1_weights[63][6] = 16'sd25;
        fc1_weights[63][7] = 16'sd53;
        fc1_weights[63][8] = 16'sd33;
        fc1_weights[63][9] = 16'sd14;
        fc1_weights[63][10] = 16'sd33;
        fc1_weights[63][11] = 16'sd30;
        fc1_weights[63][12] = 16'sd-27;
        fc1_weights[63][13] = 16'sd-45;
        fc1_weights[63][14] = 16'sd-22;
        fc1_weights[63][15] = 16'sd30;
        fc1_weights[63][16] = 16'sd-3;
        fc1_weights[63][17] = 16'sd4;
        fc1_weights[63][18] = 16'sd23;
        fc1_weights[63][19] = 16'sd-38;
        fc1_weights[63][20] = 16'sd-53;
        fc1_weights[63][21] = 16'sd-34;
        fc1_weights[63][22] = 16'sd-38;
        fc1_weights[63][23] = 16'sd-10;
        fc1_weights[63][24] = 16'sd40;
        fc1_weights[63][25] = 16'sd13;
        fc1_weights[63][26] = 16'sd16;
        fc1_weights[63][27] = 16'sd-56;
        fc1_weights[63][28] = 16'sd-62;
        fc1_weights[63][29] = 16'sd-14;
        fc1_weights[63][30] = 16'sd5;
        fc1_weights[63][31] = 16'sd20;
        fc1_weights[63][32] = 16'sd19;
        fc1_weights[63][33] = 16'sd35;
        fc1_weights[63][34] = 16'sd48;
        fc1_weights[63][35] = 16'sd56;
        fc1_weights[63][36] = 16'sd52;
        fc1_weights[63][37] = 16'sd50;
        fc1_weights[63][38] = 16'sd11;
        fc1_weights[63][39] = 16'sd-96;
        fc1_weights[63][40] = 16'sd42;
        fc1_weights[63][41] = 16'sd13;
        fc1_weights[63][42] = 16'sd-1;
        fc1_weights[63][43] = 16'sd38;
        fc1_weights[63][44] = 16'sd-6;
        fc1_weights[63][45] = 16'sd-64;
        fc1_weights[63][46] = 16'sd-22;
        fc1_weights[63][47] = 16'sd-10;
        fc1_weights[63][48] = 16'sd21;
        fc1_weights[63][49] = 16'sd40;
        fc1_weights[63][50] = 16'sd-14;
        fc1_weights[63][51] = 16'sd5;
        fc1_weights[63][52] = 16'sd-27;
        fc1_weights[63][53] = 16'sd-13;
        fc1_weights[63][54] = 16'sd-33;
        fc1_weights[63][55] = 16'sd-39;
        fc1_weights[63][56] = 16'sd-8;
        fc1_weights[63][57] = 16'sd24;
        fc1_weights[63][58] = 16'sd7;
        fc1_weights[63][59] = 16'sd-5;
        fc1_weights[63][60] = 16'sd21;
        fc1_weights[63][61] = 16'sd-5;
        fc1_weights[63][62] = 16'sd-2;
        fc1_weights[63][63] = 16'sd0;
        fc1_weights[63][64] = 16'sd3;
        fc1_weights[63][65] = 16'sd1;
        fc1_weights[63][66] = 16'sd2;
        fc1_weights[63][67] = 16'sd11;
        fc1_weights[63][68] = 16'sd12;
        fc1_weights[63][69] = 16'sd15;
        fc1_weights[63][70] = 16'sd0;
        fc1_weights[63][71] = 16'sd-44;
        fc1_weights[63][72] = 16'sd6;
        fc1_weights[63][73] = 16'sd-15;
        fc1_weights[63][74] = 16'sd-23;
        fc1_weights[63][75] = 16'sd-5;
        fc1_weights[63][76] = 16'sd32;
        fc1_weights[63][77] = 16'sd28;
        fc1_weights[63][78] = 16'sd-15;
        fc1_weights[63][79] = 16'sd-4;
        fc1_weights[63][80] = 16'sd-46;
        fc1_weights[63][81] = 16'sd0;
        fc1_weights[63][82] = 16'sd-18;
        fc1_weights[63][83] = 16'sd-14;
        fc1_weights[63][84] = 16'sd-11;
        fc1_weights[63][85] = 16'sd-44;
        fc1_weights[63][86] = 16'sd-28;
        fc1_weights[63][87] = 16'sd-19;
        fc1_weights[63][88] = 16'sd-32;
        fc1_weights[63][89] = 16'sd18;
        fc1_weights[63][90] = 16'sd-62;
        fc1_weights[63][91] = 16'sd-4;
        fc1_weights[63][92] = 16'sd-19;
        fc1_weights[63][93] = 16'sd77;
        fc1_weights[63][94] = 16'sd-18;
        fc1_weights[63][95] = 16'sd3;
        fc1_weights[63][96] = 16'sd-53;
        fc1_weights[63][97] = 16'sd-50;
        fc1_weights[63][98] = 16'sd-18;
        fc1_weights[63][99] = 16'sd-25;
        fc1_weights[63][100] = 16'sd17;
        fc1_weights[63][101] = 16'sd0;
        fc1_weights[63][102] = 16'sd18;
        fc1_weights[63][103] = 16'sd-1;
        fc1_weights[63][104] = 16'sd-29;
        fc1_weights[63][105] = 16'sd-24;
        fc1_weights[63][106] = 16'sd-38;
        fc1_weights[63][107] = 16'sd-46;
        fc1_weights[63][108] = 16'sd-34;
        fc1_weights[63][109] = 16'sd-5;
        fc1_weights[63][110] = 16'sd10;
        fc1_weights[63][111] = 16'sd-4;
        fc1_weights[63][112] = 16'sd17;
        fc1_weights[63][113] = 16'sd7;
        fc1_weights[63][114] = 16'sd55;
        fc1_weights[63][115] = 16'sd-10;
        fc1_weights[63][116] = 16'sd10;
        fc1_weights[63][117] = 16'sd32;
        fc1_weights[63][118] = 16'sd-8;
        fc1_weights[63][119] = 16'sd9;
        fc1_weights[63][120] = 16'sd-42;
        fc1_weights[63][121] = 16'sd-18;
        fc1_weights[63][122] = 16'sd-14;
        fc1_weights[63][123] = 16'sd-14;
        fc1_weights[63][124] = 16'sd-48;
        fc1_weights[63][125] = 16'sd-16;
        fc1_weights[63][126] = 16'sd-29;
        fc1_weights[63][127] = 16'sd-15;
        fc1_weights[63][128] = 16'sd-10;
        fc1_weights[63][129] = 16'sd-47;
        fc1_weights[63][130] = 16'sd-19;
        fc1_weights[63][131] = 16'sd-44;
        fc1_weights[63][132] = 16'sd0;
        fc1_weights[63][133] = 16'sd-17;
        fc1_weights[63][134] = 16'sd-2;
        fc1_weights[63][135] = 16'sd42;
        fc1_weights[63][136] = 16'sd14;
        fc1_weights[63][137] = 16'sd-7;
        fc1_weights[63][138] = 16'sd62;
        fc1_weights[63][139] = 16'sd26;
        fc1_weights[63][140] = 16'sd35;
        fc1_weights[63][141] = 16'sd-10;
        fc1_weights[63][142] = 16'sd24;
        fc1_weights[63][143] = 16'sd8;
        fc1_weights[63][144] = 16'sd71;
        fc1_weights[63][145] = 16'sd21;
        fc1_weights[63][146] = 16'sd29;
        fc1_weights[63][147] = 16'sd16;
        fc1_weights[63][148] = 16'sd0;
        fc1_weights[63][149] = 16'sd13;
        fc1_weights[63][150] = 16'sd12;
        fc1_weights[63][151] = 16'sd16;
        fc1_weights[63][152] = 16'sd13;
        fc1_weights[63][153] = 16'sd-6;
        fc1_weights[63][154] = 16'sd10;
        fc1_weights[63][155] = 16'sd16;
        fc1_weights[63][156] = 16'sd-1;
        fc1_weights[63][157] = 16'sd9;
        fc1_weights[63][158] = 16'sd-3;
        fc1_weights[63][159] = 16'sd49;
        fc1_weights[63][160] = 16'sd19;
        fc1_weights[63][161] = 16'sd-22;
        fc1_weights[63][162] = 16'sd42;
        fc1_weights[63][163] = 16'sd16;
        fc1_weights[63][164] = 16'sd35;
        fc1_weights[63][165] = 16'sd12;
        fc1_weights[63][166] = 16'sd48;
        fc1_weights[63][167] = 16'sd9;
        fc1_weights[63][168] = 16'sd67;
        fc1_weights[63][169] = 16'sd-2;
        fc1_weights[63][170] = 16'sd-9;
        fc1_weights[63][171] = 16'sd40;
        fc1_weights[63][172] = 16'sd50;
        fc1_weights[63][173] = 16'sd42;
        fc1_weights[63][174] = 16'sd25;
        fc1_weights[63][175] = 16'sd33;
        fc1_weights[63][176] = 16'sd25;
        fc1_weights[63][177] = 16'sd50;
        fc1_weights[63][178] = 16'sd-3;
        fc1_weights[63][179] = 16'sd53;
        fc1_weights[63][180] = 16'sd56;
        fc1_weights[63][181] = 16'sd5;
        fc1_weights[63][182] = 16'sd25;
        fc1_weights[63][183] = 16'sd29;
        fc1_weights[63][184] = 16'sd-19;
        fc1_weights[63][185] = 16'sd49;
        fc1_weights[63][186] = 16'sd-7;
        fc1_weights[63][187] = 16'sd9;
        fc1_weights[63][188] = 16'sd36;
        fc1_weights[63][189] = 16'sd-14;
        fc1_weights[63][190] = 16'sd7;
        fc1_weights[63][191] = 16'sd36;
        fc1_weights[63][192] = 16'sd-15;
        fc1_weights[63][193] = 16'sd-4;
        fc1_weights[63][194] = 16'sd-1;
        fc1_weights[63][195] = 16'sd-5;
        fc1_weights[63][196] = 16'sd-32;
        fc1_weights[63][197] = 16'sd29;
        fc1_weights[63][198] = 16'sd42;
        fc1_weights[63][199] = 16'sd20;
        fc1_weights[63][200] = 16'sd3;
        fc1_weights[63][201] = 16'sd22;
        fc1_weights[63][202] = 16'sd-6;
        fc1_weights[63][203] = 16'sd14;
        fc1_weights[63][204] = 16'sd38;
        fc1_weights[63][205] = 16'sd48;
        fc1_weights[63][206] = 16'sd-11;
        fc1_weights[63][207] = 16'sd-24;
        fc1_weights[64][0] = 16'sd20;
        fc1_weights[64][1] = 16'sd55;
        fc1_weights[64][2] = 16'sd-18;
        fc1_weights[64][3] = 16'sd-1;
        fc1_weights[64][4] = 16'sd13;
        fc1_weights[64][5] = 16'sd24;
        fc1_weights[64][6] = 16'sd18;
        fc1_weights[64][7] = 16'sd16;
        fc1_weights[64][8] = 16'sd-81;
        fc1_weights[64][9] = 16'sd-84;
        fc1_weights[64][10] = 16'sd-61;
        fc1_weights[64][11] = 16'sd-16;
        fc1_weights[64][12] = 16'sd41;
        fc1_weights[64][13] = 16'sd12;
        fc1_weights[64][14] = 16'sd64;
        fc1_weights[64][15] = 16'sd6;
        fc1_weights[64][16] = 16'sd10;
        fc1_weights[64][17] = 16'sd57;
        fc1_weights[64][18] = 16'sd8;
        fc1_weights[64][19] = 16'sd9;
        fc1_weights[64][20] = 16'sd-5;
        fc1_weights[64][21] = 16'sd10;
        fc1_weights[64][22] = 16'sd-32;
        fc1_weights[64][23] = 16'sd-30;
        fc1_weights[64][24] = 16'sd-19;
        fc1_weights[64][25] = 16'sd-33;
        fc1_weights[64][26] = 16'sd8;
        fc1_weights[64][27] = 16'sd-26;
        fc1_weights[64][28] = 16'sd-11;
        fc1_weights[64][29] = 16'sd42;
        fc1_weights[64][30] = 16'sd-4;
        fc1_weights[64][31] = 16'sd-2;
        fc1_weights[64][32] = 16'sd-31;
        fc1_weights[64][33] = 16'sd-1;
        fc1_weights[64][34] = 16'sd2;
        fc1_weights[64][35] = 16'sd-45;
        fc1_weights[64][36] = 16'sd-97;
        fc1_weights[64][37] = 16'sd-112;
        fc1_weights[64][38] = 16'sd-59;
        fc1_weights[64][39] = 16'sd16;
        fc1_weights[64][40] = 16'sd-38;
        fc1_weights[64][41] = 16'sd54;
        fc1_weights[64][42] = 16'sd20;
        fc1_weights[64][43] = 16'sd-28;
        fc1_weights[64][44] = 16'sd-48;
        fc1_weights[64][45] = 16'sd4;
        fc1_weights[64][46] = 16'sd-4;
        fc1_weights[64][47] = 16'sd28;
        fc1_weights[64][48] = 16'sd-29;
        fc1_weights[64][49] = 16'sd-19;
        fc1_weights[64][50] = 16'sd5;
        fc1_weights[64][51] = 16'sd50;
        fc1_weights[64][52] = 16'sd-42;
        fc1_weights[64][53] = 16'sd-38;
        fc1_weights[64][54] = 16'sd-40;
        fc1_weights[64][55] = 16'sd1;
        fc1_weights[64][56] = 16'sd13;
        fc1_weights[64][57] = 16'sd-13;
        fc1_weights[64][58] = 16'sd-3;
        fc1_weights[64][59] = 16'sd5;
        fc1_weights[64][60] = 16'sd19;
        fc1_weights[64][61] = 16'sd-7;
        fc1_weights[64][62] = 16'sd-5;
        fc1_weights[64][63] = 16'sd-31;
        fc1_weights[64][64] = 16'sd45;
        fc1_weights[64][65] = 16'sd57;
        fc1_weights[64][66] = 16'sd17;
        fc1_weights[64][67] = 16'sd22;
        fc1_weights[64][68] = 16'sd-37;
        fc1_weights[64][69] = 16'sd-22;
        fc1_weights[64][70] = 16'sd37;
        fc1_weights[64][71] = 16'sd46;
        fc1_weights[64][72] = 16'sd-3;
        fc1_weights[64][73] = 16'sd45;
        fc1_weights[64][74] = 16'sd40;
        fc1_weights[64][75] = 16'sd15;
        fc1_weights[64][76] = 16'sd1;
        fc1_weights[64][77] = 16'sd65;
        fc1_weights[64][78] = 16'sd-41;
        fc1_weights[64][79] = 16'sd-44;
        fc1_weights[64][80] = 16'sd4;
        fc1_weights[64][81] = 16'sd60;
        fc1_weights[64][82] = 16'sd-13;
        fc1_weights[64][83] = 16'sd50;
        fc1_weights[64][84] = 16'sd-26;
        fc1_weights[64][85] = 16'sd-34;
        fc1_weights[64][86] = 16'sd-8;
        fc1_weights[64][87] = 16'sd28;
        fc1_weights[64][88] = 16'sd76;
        fc1_weights[64][89] = 16'sd-91;
        fc1_weights[64][90] = 16'sd-3;
        fc1_weights[64][91] = 16'sd-4;
        fc1_weights[64][92] = 16'sd-21;
        fc1_weights[64][93] = 16'sd14;
        fc1_weights[64][94] = 16'sd-28;
        fc1_weights[64][95] = 16'sd14;
        fc1_weights[64][96] = 16'sd33;
        fc1_weights[64][97] = 16'sd45;
        fc1_weights[64][98] = 16'sd44;
        fc1_weights[64][99] = 16'sd-20;
        fc1_weights[64][100] = 16'sd22;
        fc1_weights[64][101] = 16'sd-5;
        fc1_weights[64][102] = 16'sd-2;
        fc1_weights[64][103] = 16'sd51;
        fc1_weights[64][104] = 16'sd28;
        fc1_weights[64][105] = 16'sd-29;
        fc1_weights[64][106] = 16'sd35;
        fc1_weights[64][107] = 16'sd56;
        fc1_weights[64][108] = 16'sd31;
        fc1_weights[64][109] = 16'sd15;
        fc1_weights[64][110] = 16'sd-37;
        fc1_weights[64][111] = 16'sd-67;
        fc1_weights[64][112] = 16'sd-37;
        fc1_weights[64][113] = 16'sd-29;
        fc1_weights[64][114] = 16'sd-14;
        fc1_weights[64][115] = 16'sd-42;
        fc1_weights[64][116] = 16'sd-41;
        fc1_weights[64][117] = 16'sd-39;
        fc1_weights[64][118] = 16'sd-12;
        fc1_weights[64][119] = 16'sd-15;
        fc1_weights[64][120] = 16'sd15;
        fc1_weights[64][121] = 16'sd-7;
        fc1_weights[64][122] = 16'sd-27;
        fc1_weights[64][123] = 16'sd-55;
        fc1_weights[64][124] = 16'sd-17;
        fc1_weights[64][125] = 16'sd-53;
        fc1_weights[64][126] = 16'sd60;
        fc1_weights[64][127] = 16'sd0;
        fc1_weights[64][128] = 16'sd20;
        fc1_weights[64][129] = 16'sd49;
        fc1_weights[64][130] = 16'sd10;
        fc1_weights[64][131] = 16'sd48;
        fc1_weights[64][132] = 16'sd18;
        fc1_weights[64][133] = 16'sd50;
        fc1_weights[64][134] = 16'sd20;
        fc1_weights[64][135] = 16'sd47;
        fc1_weights[64][136] = 16'sd27;
        fc1_weights[64][137] = 16'sd-36;
        fc1_weights[64][138] = 16'sd43;
        fc1_weights[64][139] = 16'sd-98;
        fc1_weights[64][140] = 16'sd-57;
        fc1_weights[64][141] = 16'sd2;
        fc1_weights[64][142] = 16'sd-44;
        fc1_weights[64][143] = 16'sd-50;
        fc1_weights[64][144] = 16'sd44;
        fc1_weights[64][145] = 16'sd24;
        fc1_weights[64][146] = 16'sd17;
        fc1_weights[64][147] = 16'sd-29;
        fc1_weights[64][148] = 16'sd-39;
        fc1_weights[64][149] = 16'sd13;
        fc1_weights[64][150] = 16'sd31;
        fc1_weights[64][151] = 16'sd91;
        fc1_weights[64][152] = 16'sd-2;
        fc1_weights[64][153] = 16'sd-38;
        fc1_weights[64][154] = 16'sd-14;
        fc1_weights[64][155] = 16'sd21;
        fc1_weights[64][156] = 16'sd-36;
        fc1_weights[64][157] = 16'sd-32;
        fc1_weights[64][158] = 16'sd-7;
        fc1_weights[64][159] = 16'sd71;
        fc1_weights[64][160] = 16'sd32;
        fc1_weights[64][161] = 16'sd57;
        fc1_weights[64][162] = 16'sd52;
        fc1_weights[64][163] = 16'sd-17;
        fc1_weights[64][164] = 16'sd-19;
        fc1_weights[64][165] = 16'sd-38;
        fc1_weights[64][166] = 16'sd-76;
        fc1_weights[64][167] = 16'sd-51;
        fc1_weights[64][168] = 16'sd-24;
        fc1_weights[64][169] = 16'sd-7;
        fc1_weights[64][170] = 16'sd6;
        fc1_weights[64][171] = 16'sd-35;
        fc1_weights[64][172] = 16'sd-31;
        fc1_weights[64][173] = 16'sd-45;
        fc1_weights[64][174] = 16'sd1;
        fc1_weights[64][175] = 16'sd-22;
        fc1_weights[64][176] = 16'sd-19;
        fc1_weights[64][177] = 16'sd41;
        fc1_weights[64][178] = 16'sd78;
        fc1_weights[64][179] = 16'sd33;
        fc1_weights[64][180] = 16'sd70;
        fc1_weights[64][181] = 16'sd68;
        fc1_weights[64][182] = 16'sd1;
        fc1_weights[64][183] = 16'sd30;
        fc1_weights[64][184] = 16'sd78;
        fc1_weights[64][185] = 16'sd29;
        fc1_weights[64][186] = 16'sd6;
        fc1_weights[64][187] = 16'sd-29;
        fc1_weights[64][188] = 16'sd-39;
        fc1_weights[64][189] = 16'sd0;
        fc1_weights[64][190] = 16'sd-2;
        fc1_weights[64][191] = 16'sd-51;
        fc1_weights[64][192] = 16'sd3;
        fc1_weights[64][193] = 16'sd-4;
        fc1_weights[64][194] = 16'sd9;
        fc1_weights[64][195] = 16'sd19;
        fc1_weights[64][196] = 16'sd48;
        fc1_weights[64][197] = 16'sd56;
        fc1_weights[64][198] = 16'sd31;
        fc1_weights[64][199] = 16'sd-19;
        fc1_weights[64][200] = 16'sd42;
        fc1_weights[64][201] = 16'sd-17;
        fc1_weights[64][202] = 16'sd8;
        fc1_weights[64][203] = 16'sd11;
        fc1_weights[64][204] = 16'sd-10;
        fc1_weights[64][205] = 16'sd7;
        fc1_weights[64][206] = 16'sd38;
        fc1_weights[64][207] = 16'sd105;
        fc1_weights[65][0] = 16'sd-8;
        fc1_weights[65][1] = 16'sd15;
        fc1_weights[65][2] = 16'sd29;
        fc1_weights[65][3] = 16'sd-15;
        fc1_weights[65][4] = 16'sd-13;
        fc1_weights[65][5] = 16'sd14;
        fc1_weights[65][6] = 16'sd33;
        fc1_weights[65][7] = 16'sd22;
        fc1_weights[65][8] = 16'sd62;
        fc1_weights[65][9] = 16'sd-8;
        fc1_weights[65][10] = 16'sd-16;
        fc1_weights[65][11] = 16'sd-81;
        fc1_weights[65][12] = 16'sd-88;
        fc1_weights[65][13] = 16'sd-32;
        fc1_weights[65][14] = 16'sd37;
        fc1_weights[65][15] = 16'sd99;
        fc1_weights[65][16] = 16'sd70;
        fc1_weights[65][17] = 16'sd18;
        fc1_weights[65][18] = 16'sd59;
        fc1_weights[65][19] = 16'sd-9;
        fc1_weights[65][20] = 16'sd23;
        fc1_weights[65][21] = 16'sd-28;
        fc1_weights[65][22] = 16'sd47;
        fc1_weights[65][23] = 16'sd-18;
        fc1_weights[65][24] = 16'sd85;
        fc1_weights[65][25] = 16'sd51;
        fc1_weights[65][26] = 16'sd42;
        fc1_weights[65][27] = 16'sd25;
        fc1_weights[65][28] = 16'sd12;
        fc1_weights[65][29] = 16'sd13;
        fc1_weights[65][30] = 16'sd33;
        fc1_weights[65][31] = 16'sd24;
        fc1_weights[65][32] = 16'sd34;
        fc1_weights[65][33] = 16'sd67;
        fc1_weights[65][34] = 16'sd22;
        fc1_weights[65][35] = 16'sd40;
        fc1_weights[65][36] = 16'sd-8;
        fc1_weights[65][37] = 16'sd-85;
        fc1_weights[65][38] = 16'sd-51;
        fc1_weights[65][39] = 16'sd-41;
        fc1_weights[65][40] = 16'sd95;
        fc1_weights[65][41] = 16'sd126;
        fc1_weights[65][42] = 16'sd-5;
        fc1_weights[65][43] = 16'sd89;
        fc1_weights[65][44] = 16'sd0;
        fc1_weights[65][45] = 16'sd-33;
        fc1_weights[65][46] = 16'sd16;
        fc1_weights[65][47] = 16'sd-37;
        fc1_weights[65][48] = 16'sd-68;
        fc1_weights[65][49] = 16'sd-7;
        fc1_weights[65][50] = 16'sd-20;
        fc1_weights[65][51] = 16'sd-30;
        fc1_weights[65][52] = 16'sd2;
        fc1_weights[65][53] = 16'sd24;
        fc1_weights[65][54] = 16'sd-31;
        fc1_weights[65][55] = 16'sd-21;
        fc1_weights[65][56] = 16'sd-16;
        fc1_weights[65][57] = 16'sd18;
        fc1_weights[65][58] = 16'sd33;
        fc1_weights[65][59] = 16'sd9;
        fc1_weights[65][60] = 16'sd-22;
        fc1_weights[65][61] = 16'sd-13;
        fc1_weights[65][62] = 16'sd-53;
        fc1_weights[65][63] = 16'sd19;
        fc1_weights[65][64] = 16'sd-61;
        fc1_weights[65][65] = 16'sd-31;
        fc1_weights[65][66] = 16'sd59;
        fc1_weights[65][67] = 16'sd63;
        fc1_weights[65][68] = 16'sd46;
        fc1_weights[65][69] = 16'sd-9;
        fc1_weights[65][70] = 16'sd18;
        fc1_weights[65][71] = 16'sd24;
        fc1_weights[65][72] = 16'sd76;
        fc1_weights[65][73] = 16'sd-25;
        fc1_weights[65][74] = 16'sd-28;
        fc1_weights[65][75] = 16'sd-67;
        fc1_weights[65][76] = 16'sd32;
        fc1_weights[65][77] = 16'sd-1;
        fc1_weights[65][78] = 16'sd-10;
        fc1_weights[65][79] = 16'sd48;
        fc1_weights[65][80] = 16'sd-5;
        fc1_weights[65][81] = 16'sd-25;
        fc1_weights[65][82] = 16'sd-32;
        fc1_weights[65][83] = 16'sd9;
        fc1_weights[65][84] = 16'sd20;
        fc1_weights[65][85] = 16'sd2;
        fc1_weights[65][86] = 16'sd3;
        fc1_weights[65][87] = 16'sd-18;
        fc1_weights[65][88] = 16'sd-97;
        fc1_weights[65][89] = 16'sd-58;
        fc1_weights[65][90] = 16'sd-23;
        fc1_weights[65][91] = 16'sd1;
        fc1_weights[65][92] = 16'sd-29;
        fc1_weights[65][93] = 16'sd44;
        fc1_weights[65][94] = 16'sd-10;
        fc1_weights[65][95] = 16'sd18;
        fc1_weights[65][96] = 16'sd-23;
        fc1_weights[65][97] = 16'sd-6;
        fc1_weights[65][98] = 16'sd85;
        fc1_weights[65][99] = 16'sd22;
        fc1_weights[65][100] = 16'sd-61;
        fc1_weights[65][101] = 16'sd-62;
        fc1_weights[65][102] = 16'sd-24;
        fc1_weights[65][103] = 16'sd-15;
        fc1_weights[65][104] = 16'sd19;
        fc1_weights[65][105] = 16'sd10;
        fc1_weights[65][106] = 16'sd26;
        fc1_weights[65][107] = 16'sd18;
        fc1_weights[65][108] = 16'sd28;
        fc1_weights[65][109] = 16'sd14;
        fc1_weights[65][110] = 16'sd16;
        fc1_weights[65][111] = 16'sd-72;
        fc1_weights[65][112] = 16'sd2;
        fc1_weights[65][113] = 16'sd1;
        fc1_weights[65][114] = 16'sd-40;
        fc1_weights[65][115] = 16'sd-16;
        fc1_weights[65][116] = 16'sd-29;
        fc1_weights[65][117] = 16'sd-17;
        fc1_weights[65][118] = 16'sd-54;
        fc1_weights[65][119] = 16'sd-26;
        fc1_weights[65][120] = 16'sd-21;
        fc1_weights[65][121] = 16'sd-27;
        fc1_weights[65][122] = 16'sd-60;
        fc1_weights[65][123] = 16'sd-43;
        fc1_weights[65][124] = 16'sd-90;
        fc1_weights[65][125] = 16'sd-39;
        fc1_weights[65][126] = 16'sd-110;
        fc1_weights[65][127] = 16'sd-61;
        fc1_weights[65][128] = 16'sd-95;
        fc1_weights[65][129] = 16'sd-65;
        fc1_weights[65][130] = 16'sd-73;
        fc1_weights[65][131] = 16'sd-33;
        fc1_weights[65][132] = 16'sd-14;
        fc1_weights[65][133] = 16'sd-24;
        fc1_weights[65][134] = 16'sd13;
        fc1_weights[65][135] = 16'sd53;
        fc1_weights[65][136] = 16'sd2;
        fc1_weights[65][137] = 16'sd-21;
        fc1_weights[65][138] = 16'sd13;
        fc1_weights[65][139] = 16'sd-34;
        fc1_weights[65][140] = 16'sd52;
        fc1_weights[65][141] = 16'sd-32;
        fc1_weights[65][142] = 16'sd50;
        fc1_weights[65][143] = 16'sd53;
        fc1_weights[65][144] = 16'sd30;
        fc1_weights[65][145] = 16'sd-33;
        fc1_weights[65][146] = 16'sd-47;
        fc1_weights[65][147] = 16'sd46;
        fc1_weights[65][148] = 16'sd-69;
        fc1_weights[65][149] = 16'sd-69;
        fc1_weights[65][150] = 16'sd-60;
        fc1_weights[65][151] = 16'sd-21;
        fc1_weights[65][152] = 16'sd15;
        fc1_weights[65][153] = 16'sd-24;
        fc1_weights[65][154] = 16'sd-20;
        fc1_weights[65][155] = 16'sd55;
        fc1_weights[65][156] = 16'sd26;
        fc1_weights[65][157] = 16'sd21;
        fc1_weights[65][158] = 16'sd66;
        fc1_weights[65][159] = 16'sd-18;
        fc1_weights[65][160] = 16'sd-45;
        fc1_weights[65][161] = 16'sd-22;
        fc1_weights[65][162] = 16'sd-58;
        fc1_weights[65][163] = 16'sd-41;
        fc1_weights[65][164] = 16'sd-44;
        fc1_weights[65][165] = 16'sd46;
        fc1_weights[65][166] = 16'sd48;
        fc1_weights[65][167] = 16'sd25;
        fc1_weights[65][168] = 16'sd-2;
        fc1_weights[65][169] = 16'sd29;
        fc1_weights[65][170] = 16'sd41;
        fc1_weights[65][171] = 16'sd15;
        fc1_weights[65][172] = 16'sd40;
        fc1_weights[65][173] = 16'sd40;
        fc1_weights[65][174] = 16'sd60;
        fc1_weights[65][175] = 16'sd27;
        fc1_weights[65][176] = 16'sd49;
        fc1_weights[65][177] = 16'sd7;
        fc1_weights[65][178] = 16'sd6;
        fc1_weights[65][179] = 16'sd27;
        fc1_weights[65][180] = 16'sd-1;
        fc1_weights[65][181] = 16'sd-11;
        fc1_weights[65][182] = 16'sd-11;
        fc1_weights[65][183] = 16'sd60;
        fc1_weights[65][184] = 16'sd11;
        fc1_weights[65][185] = 16'sd-15;
        fc1_weights[65][186] = 16'sd-10;
        fc1_weights[65][187] = 16'sd-67;
        fc1_weights[65][188] = 16'sd-66;
        fc1_weights[65][189] = 16'sd-38;
        fc1_weights[65][190] = 16'sd63;
        fc1_weights[65][191] = 16'sd27;
        fc1_weights[65][192] = 16'sd2;
        fc1_weights[65][193] = 16'sd6;
        fc1_weights[65][194] = 16'sd-10;
        fc1_weights[65][195] = 16'sd-2;
        fc1_weights[65][196] = 16'sd10;
        fc1_weights[65][197] = 16'sd16;
        fc1_weights[65][198] = 16'sd11;
        fc1_weights[65][199] = 16'sd39;
        fc1_weights[65][200] = 16'sd-15;
        fc1_weights[65][201] = 16'sd-53;
        fc1_weights[65][202] = 16'sd-5;
        fc1_weights[65][203] = 16'sd57;
        fc1_weights[65][204] = 16'sd-1;
        fc1_weights[65][205] = 16'sd2;
        fc1_weights[65][206] = 16'sd-58;
        fc1_weights[65][207] = 16'sd-7;
        fc1_weights[66][0] = 16'sd5;
        fc1_weights[66][1] = 16'sd30;
        fc1_weights[66][2] = 16'sd-18;
        fc1_weights[66][3] = 16'sd-15;
        fc1_weights[66][4] = 16'sd-40;
        fc1_weights[66][5] = 16'sd-28;
        fc1_weights[66][6] = 16'sd-10;
        fc1_weights[66][7] = 16'sd55;
        fc1_weights[66][8] = 16'sd33;
        fc1_weights[66][9] = 16'sd23;
        fc1_weights[66][10] = 16'sd53;
        fc1_weights[66][11] = 16'sd57;
        fc1_weights[66][12] = 16'sd-25;
        fc1_weights[66][13] = 16'sd-94;
        fc1_weights[66][14] = 16'sd-56;
        fc1_weights[66][15] = 16'sd5;
        fc1_weights[66][16] = 16'sd12;
        fc1_weights[66][17] = 16'sd27;
        fc1_weights[66][18] = 16'sd28;
        fc1_weights[66][19] = 16'sd-45;
        fc1_weights[66][20] = 16'sd25;
        fc1_weights[66][21] = 16'sd-50;
        fc1_weights[66][22] = 16'sd-41;
        fc1_weights[66][23] = 16'sd-44;
        fc1_weights[66][24] = 16'sd11;
        fc1_weights[66][25] = 16'sd0;
        fc1_weights[66][26] = 16'sd18;
        fc1_weights[66][27] = 16'sd-29;
        fc1_weights[66][28] = 16'sd-23;
        fc1_weights[66][29] = 16'sd48;
        fc1_weights[66][30] = 16'sd27;
        fc1_weights[66][31] = 16'sd20;
        fc1_weights[66][32] = 16'sd68;
        fc1_weights[66][33] = 16'sd-68;
        fc1_weights[66][34] = 16'sd86;
        fc1_weights[66][35] = 16'sd52;
        fc1_weights[66][36] = 16'sd15;
        fc1_weights[66][37] = 16'sd110;
        fc1_weights[66][38] = 16'sd61;
        fc1_weights[66][39] = 16'sd-86;
        fc1_weights[66][40] = 16'sd59;
        fc1_weights[66][41] = 16'sd-8;
        fc1_weights[66][42] = 16'sd-8;
        fc1_weights[66][43] = 16'sd22;
        fc1_weights[66][44] = 16'sd-18;
        fc1_weights[66][45] = 16'sd-15;
        fc1_weights[66][46] = 16'sd0;
        fc1_weights[66][47] = 16'sd-75;
        fc1_weights[66][48] = 16'sd21;
        fc1_weights[66][49] = 16'sd31;
        fc1_weights[66][50] = 16'sd-26;
        fc1_weights[66][51] = 16'sd6;
        fc1_weights[66][52] = 16'sd-64;
        fc1_weights[66][53] = 16'sd-67;
        fc1_weights[66][54] = 16'sd-5;
        fc1_weights[66][55] = 16'sd14;
        fc1_weights[66][56] = 16'sd21;
        fc1_weights[66][57] = 16'sd37;
        fc1_weights[66][58] = 16'sd-31;
        fc1_weights[66][59] = 16'sd-53;
        fc1_weights[66][60] = 16'sd50;
        fc1_weights[66][61] = 16'sd11;
        fc1_weights[66][62] = 16'sd2;
        fc1_weights[66][63] = 16'sd81;
        fc1_weights[66][64] = 16'sd102;
        fc1_weights[66][65] = 16'sd-36;
        fc1_weights[66][66] = 16'sd13;
        fc1_weights[66][67] = 16'sd-51;
        fc1_weights[66][68] = 16'sd-4;
        fc1_weights[66][69] = 16'sd-6;
        fc1_weights[66][70] = 16'sd31;
        fc1_weights[66][71] = 16'sd-23;
        fc1_weights[66][72] = 16'sd-22;
        fc1_weights[66][73] = 16'sd-10;
        fc1_weights[66][74] = 16'sd48;
        fc1_weights[66][75] = 16'sd-43;
        fc1_weights[66][76] = 16'sd32;
        fc1_weights[66][77] = 16'sd72;
        fc1_weights[66][78] = 16'sd19;
        fc1_weights[66][79] = 16'sd33;
        fc1_weights[66][80] = 16'sd-9;
        fc1_weights[66][81] = 16'sd-58;
        fc1_weights[66][82] = 16'sd-39;
        fc1_weights[66][83] = 16'sd-32;
        fc1_weights[66][84] = 16'sd-36;
        fc1_weights[66][85] = 16'sd-121;
        fc1_weights[66][86] = 16'sd-43;
        fc1_weights[66][87] = 16'sd57;
        fc1_weights[66][88] = 16'sd-13;
        fc1_weights[66][89] = 16'sd28;
        fc1_weights[66][90] = 16'sd79;
        fc1_weights[66][91] = 16'sd-4;
        fc1_weights[66][92] = 16'sd13;
        fc1_weights[66][93] = 16'sd3;
        fc1_weights[66][94] = 16'sd-44;
        fc1_weights[66][95] = 16'sd53;
        fc1_weights[66][96] = 16'sd-34;
        fc1_weights[66][97] = 16'sd42;
        fc1_weights[66][98] = 16'sd1;
        fc1_weights[66][99] = 16'sd-25;
        fc1_weights[66][100] = 16'sd31;
        fc1_weights[66][101] = 16'sd26;
        fc1_weights[66][102] = 16'sd-17;
        fc1_weights[66][103] = 16'sd25;
        fc1_weights[66][104] = 16'sd-33;
        fc1_weights[66][105] = 16'sd-25;
        fc1_weights[66][106] = 16'sd-46;
        fc1_weights[66][107] = 16'sd-68;
        fc1_weights[66][108] = 16'sd-14;
        fc1_weights[66][109] = 16'sd-25;
        fc1_weights[66][110] = 16'sd-54;
        fc1_weights[66][111] = 16'sd-52;
        fc1_weights[66][112] = 16'sd35;
        fc1_weights[66][113] = 16'sd45;
        fc1_weights[66][114] = 16'sd26;
        fc1_weights[66][115] = 16'sd70;
        fc1_weights[66][116] = 16'sd46;
        fc1_weights[66][117] = 16'sd84;
        fc1_weights[66][118] = 16'sd-4;
        fc1_weights[66][119] = 16'sd13;
        fc1_weights[66][120] = 16'sd-9;
        fc1_weights[66][121] = 16'sd1;
        fc1_weights[66][122] = 16'sd20;
        fc1_weights[66][123] = 16'sd84;
        fc1_weights[66][124] = 16'sd-50;
        fc1_weights[66][125] = 16'sd-35;
        fc1_weights[66][126] = 16'sd21;
        fc1_weights[66][127] = 16'sd-5;
        fc1_weights[66][128] = 16'sd7;
        fc1_weights[66][129] = 16'sd40;
        fc1_weights[66][130] = 16'sd-77;
        fc1_weights[66][131] = 16'sd-37;
        fc1_weights[66][132] = 16'sd13;
        fc1_weights[66][133] = 16'sd-58;
        fc1_weights[66][134] = 16'sd-27;
        fc1_weights[66][135] = 16'sd-31;
        fc1_weights[66][136] = 16'sd-41;
        fc1_weights[66][137] = 16'sd-48;
        fc1_weights[66][138] = 16'sd101;
        fc1_weights[66][139] = 16'sd9;
        fc1_weights[66][140] = 16'sd-10;
        fc1_weights[66][141] = 16'sd-68;
        fc1_weights[66][142] = 16'sd17;
        fc1_weights[66][143] = 16'sd19;
        fc1_weights[66][144] = 16'sd92;
        fc1_weights[66][145] = 16'sd-9;
        fc1_weights[66][146] = 16'sd11;
        fc1_weights[66][147] = 16'sd-23;
        fc1_weights[66][148] = 16'sd22;
        fc1_weights[66][149] = 16'sd26;
        fc1_weights[66][150] = 16'sd9;
        fc1_weights[66][151] = 16'sd76;
        fc1_weights[66][152] = 16'sd-36;
        fc1_weights[66][153] = 16'sd14;
        fc1_weights[66][154] = 16'sd22;
        fc1_weights[66][155] = 16'sd47;
        fc1_weights[66][156] = 16'sd-7;
        fc1_weights[66][157] = 16'sd-27;
        fc1_weights[66][158] = 16'sd-17;
        fc1_weights[66][159] = 16'sd-4;
        fc1_weights[66][160] = 16'sd-25;
        fc1_weights[66][161] = 16'sd-78;
        fc1_weights[66][162] = 16'sd64;
        fc1_weights[66][163] = 16'sd-24;
        fc1_weights[66][164] = 16'sd-19;
        fc1_weights[66][165] = 16'sd-22;
        fc1_weights[66][166] = 16'sd-2;
        fc1_weights[66][167] = 16'sd-4;
        fc1_weights[66][168] = 16'sd58;
        fc1_weights[66][169] = 16'sd7;
        fc1_weights[66][170] = 16'sd66;
        fc1_weights[66][171] = 16'sd26;
        fc1_weights[66][172] = 16'sd35;
        fc1_weights[66][173] = 16'sd-17;
        fc1_weights[66][174] = 16'sd-24;
        fc1_weights[66][175] = 16'sd-27;
        fc1_weights[66][176] = 16'sd6;
        fc1_weights[66][177] = 16'sd101;
        fc1_weights[66][178] = 16'sd-16;
        fc1_weights[66][179] = 16'sd40;
        fc1_weights[66][180] = 16'sd81;
        fc1_weights[66][181] = 16'sd-4;
        fc1_weights[66][182] = 16'sd40;
        fc1_weights[66][183] = 16'sd-7;
        fc1_weights[66][184] = 16'sd-18;
        fc1_weights[66][185] = 16'sd79;
        fc1_weights[66][186] = 16'sd-29;
        fc1_weights[66][187] = 16'sd-10;
        fc1_weights[66][188] = 16'sd50;
        fc1_weights[66][189] = 16'sd-87;
        fc1_weights[66][190] = 16'sd31;
        fc1_weights[66][191] = 16'sd40;
        fc1_weights[66][192] = 16'sd-30;
        fc1_weights[66][193] = 16'sd-15;
        fc1_weights[66][194] = 16'sd25;
        fc1_weights[66][195] = 16'sd45;
        fc1_weights[66][196] = 16'sd-28;
        fc1_weights[66][197] = 16'sd66;
        fc1_weights[66][198] = 16'sd-4;
        fc1_weights[66][199] = 16'sd-52;
        fc1_weights[66][200] = 16'sd26;
        fc1_weights[66][201] = 16'sd-46;
        fc1_weights[66][202] = 16'sd-37;
        fc1_weights[66][203] = 16'sd9;
        fc1_weights[66][204] = 16'sd21;
        fc1_weights[66][205] = 16'sd25;
        fc1_weights[66][206] = 16'sd-8;
        fc1_weights[66][207] = 16'sd16;
        fc1_weights[67][0] = 16'sd-34;
        fc1_weights[67][1] = 16'sd-18;
        fc1_weights[67][2] = 16'sd-36;
        fc1_weights[67][3] = 16'sd-12;
        fc1_weights[67][4] = 16'sd-30;
        fc1_weights[67][5] = 16'sd16;
        fc1_weights[67][6] = 16'sd10;
        fc1_weights[67][7] = 16'sd33;
        fc1_weights[67][8] = 16'sd9;
        fc1_weights[67][9] = 16'sd-18;
        fc1_weights[67][10] = 16'sd14;
        fc1_weights[67][11] = 16'sd9;
        fc1_weights[67][12] = 16'sd45;
        fc1_weights[67][13] = 16'sd63;
        fc1_weights[67][14] = 16'sd24;
        fc1_weights[67][15] = 16'sd-50;
        fc1_weights[67][16] = 16'sd7;
        fc1_weights[67][17] = 16'sd14;
        fc1_weights[67][18] = 16'sd-7;
        fc1_weights[67][19] = 16'sd4;
        fc1_weights[67][20] = 16'sd-9;
        fc1_weights[67][21] = 16'sd14;
        fc1_weights[67][22] = 16'sd23;
        fc1_weights[67][23] = 16'sd10;
        fc1_weights[67][24] = 16'sd-9;
        fc1_weights[67][25] = 16'sd0;
        fc1_weights[67][26] = 16'sd-23;
        fc1_weights[67][27] = 16'sd-72;
        fc1_weights[67][28] = 16'sd0;
        fc1_weights[67][29] = 16'sd-26;
        fc1_weights[67][30] = 16'sd-46;
        fc1_weights[67][31] = 16'sd3;
        fc1_weights[67][32] = 16'sd6;
        fc1_weights[67][33] = 16'sd53;
        fc1_weights[67][34] = 16'sd-5;
        fc1_weights[67][35] = 16'sd-27;
        fc1_weights[67][36] = 16'sd0;
        fc1_weights[67][37] = 16'sd-3;
        fc1_weights[67][38] = 16'sd9;
        fc1_weights[67][39] = 16'sd36;
        fc1_weights[67][40] = 16'sd-23;
        fc1_weights[67][41] = 16'sd-57;
        fc1_weights[67][42] = 16'sd-20;
        fc1_weights[67][43] = 16'sd-47;
        fc1_weights[67][44] = 16'sd-14;
        fc1_weights[67][45] = 16'sd13;
        fc1_weights[67][46] = 16'sd-7;
        fc1_weights[67][47] = 16'sd46;
        fc1_weights[67][48] = 16'sd-12;
        fc1_weights[67][49] = 16'sd6;
        fc1_weights[67][50] = 16'sd-2;
        fc1_weights[67][51] = 16'sd4;
        fc1_weights[67][52] = 16'sd-8;
        fc1_weights[67][53] = 16'sd-20;
        fc1_weights[67][54] = 16'sd-18;
        fc1_weights[67][55] = 16'sd6;
        fc1_weights[67][56] = 16'sd-34;
        fc1_weights[67][57] = 16'sd-37;
        fc1_weights[67][58] = 16'sd-25;
        fc1_weights[67][59] = 16'sd-8;
        fc1_weights[67][60] = 16'sd-46;
        fc1_weights[67][61] = 16'sd-65;
        fc1_weights[67][62] = 16'sd7;
        fc1_weights[67][63] = 16'sd15;
        fc1_weights[67][64] = 16'sd-9;
        fc1_weights[67][65] = 16'sd44;
        fc1_weights[67][66] = 16'sd53;
        fc1_weights[67][67] = 16'sd-1;
        fc1_weights[67][68] = 16'sd32;
        fc1_weights[67][69] = 16'sd1;
        fc1_weights[67][70] = 16'sd43;
        fc1_weights[67][71] = 16'sd40;
        fc1_weights[67][72] = 16'sd31;
        fc1_weights[67][73] = 16'sd49;
        fc1_weights[67][74] = 16'sd17;
        fc1_weights[67][75] = 16'sd37;
        fc1_weights[67][76] = 16'sd-28;
        fc1_weights[67][77] = 16'sd17;
        fc1_weights[67][78] = 16'sd-36;
        fc1_weights[67][79] = 16'sd13;
        fc1_weights[67][80] = 16'sd-10;
        fc1_weights[67][81] = 16'sd-5;
        fc1_weights[67][82] = 16'sd-43;
        fc1_weights[67][83] = 16'sd22;
        fc1_weights[67][84] = 16'sd-5;
        fc1_weights[67][85] = 16'sd4;
        fc1_weights[67][86] = 16'sd6;
        fc1_weights[67][87] = 16'sd-56;
        fc1_weights[67][88] = 16'sd16;
        fc1_weights[67][89] = 16'sd-29;
        fc1_weights[67][90] = 16'sd-15;
        fc1_weights[67][91] = 16'sd-6;
        fc1_weights[67][92] = 16'sd-6;
        fc1_weights[67][93] = 16'sd-15;
        fc1_weights[67][94] = 16'sd-27;
        fc1_weights[67][95] = 16'sd12;
        fc1_weights[67][96] = 16'sd41;
        fc1_weights[67][97] = 16'sd-15;
        fc1_weights[67][98] = 16'sd26;
        fc1_weights[67][99] = 16'sd44;
        fc1_weights[67][100] = 16'sd18;
        fc1_weights[67][101] = 16'sd50;
        fc1_weights[67][102] = 16'sd40;
        fc1_weights[67][103] = 16'sd8;
        fc1_weights[67][104] = 16'sd-14;
        fc1_weights[67][105] = 16'sd-25;
        fc1_weights[67][106] = 16'sd-3;
        fc1_weights[67][107] = 16'sd-26;
        fc1_weights[67][108] = 16'sd-6;
        fc1_weights[67][109] = 16'sd8;
        fc1_weights[67][110] = 16'sd-11;
        fc1_weights[67][111] = 16'sd-12;
        fc1_weights[67][112] = 16'sd-9;
        fc1_weights[67][113] = 16'sd-87;
        fc1_weights[67][114] = 16'sd-17;
        fc1_weights[67][115] = 16'sd-24;
        fc1_weights[67][116] = 16'sd-2;
        fc1_weights[67][117] = 16'sd-12;
        fc1_weights[67][118] = 16'sd-20;
        fc1_weights[67][119] = 16'sd2;
        fc1_weights[67][120] = 16'sd13;
        fc1_weights[67][121] = 16'sd10;
        fc1_weights[67][122] = 16'sd9;
        fc1_weights[67][123] = 16'sd0;
        fc1_weights[67][124] = 16'sd17;
        fc1_weights[67][125] = 16'sd3;
        fc1_weights[67][126] = 16'sd3;
        fc1_weights[67][127] = 16'sd-48;
        fc1_weights[67][128] = 16'sd-18;
        fc1_weights[67][129] = 16'sd5;
        fc1_weights[67][130] = 16'sd2;
        fc1_weights[67][131] = 16'sd46;
        fc1_weights[67][132] = 16'sd41;
        fc1_weights[67][133] = 16'sd12;
        fc1_weights[67][134] = 16'sd11;
        fc1_weights[67][135] = 16'sd-20;
        fc1_weights[67][136] = 16'sd-32;
        fc1_weights[67][137] = 16'sd27;
        fc1_weights[67][138] = 16'sd-17;
        fc1_weights[67][139] = 16'sd-14;
        fc1_weights[67][140] = 16'sd17;
        fc1_weights[67][141] = 16'sd46;
        fc1_weights[67][142] = 16'sd-29;
        fc1_weights[67][143] = 16'sd-40;
        fc1_weights[67][144] = 16'sd-40;
        fc1_weights[67][145] = 16'sd-32;
        fc1_weights[67][146] = 16'sd-49;
        fc1_weights[67][147] = 16'sd5;
        fc1_weights[67][148] = 16'sd-17;
        fc1_weights[67][149] = 16'sd-18;
        fc1_weights[67][150] = 16'sd6;
        fc1_weights[67][151] = 16'sd11;
        fc1_weights[67][152] = 16'sd0;
        fc1_weights[67][153] = 16'sd-9;
        fc1_weights[67][154] = 16'sd21;
        fc1_weights[67][155] = 16'sd-34;
        fc1_weights[67][156] = 16'sd29;
        fc1_weights[67][157] = 16'sd38;
        fc1_weights[67][158] = 16'sd2;
        fc1_weights[67][159] = 16'sd22;
        fc1_weights[67][160] = 16'sd33;
        fc1_weights[67][161] = 16'sd49;
        fc1_weights[67][162] = 16'sd-15;
        fc1_weights[67][163] = 16'sd-13;
        fc1_weights[67][164] = 16'sd12;
        fc1_weights[67][165] = 16'sd24;
        fc1_weights[67][166] = 16'sd5;
        fc1_weights[67][167] = 16'sd-23;
        fc1_weights[67][168] = 16'sd-26;
        fc1_weights[67][169] = 16'sd-22;
        fc1_weights[67][170] = 16'sd-18;
        fc1_weights[67][171] = 16'sd-53;
        fc1_weights[67][172] = 16'sd-29;
        fc1_weights[67][173] = 16'sd-2;
        fc1_weights[67][174] = 16'sd21;
        fc1_weights[67][175] = 16'sd14;
        fc1_weights[67][176] = 16'sd23;
        fc1_weights[67][177] = 16'sd0;
        fc1_weights[67][178] = 16'sd3;
        fc1_weights[67][179] = 16'sd-21;
        fc1_weights[67][180] = 16'sd11;
        fc1_weights[67][181] = 16'sd-18;
        fc1_weights[67][182] = 16'sd50;
        fc1_weights[67][183] = 16'sd2;
        fc1_weights[67][184] = 16'sd18;
        fc1_weights[67][185] = 16'sd-39;
        fc1_weights[67][186] = 16'sd-29;
        fc1_weights[67][187] = 16'sd-42;
        fc1_weights[67][188] = 16'sd-22;
        fc1_weights[67][189] = 16'sd-36;
        fc1_weights[67][190] = 16'sd-31;
        fc1_weights[67][191] = 16'sd-33;
        fc1_weights[67][192] = 16'sd-21;
        fc1_weights[67][193] = 16'sd-38;
        fc1_weights[67][194] = 16'sd-4;
        fc1_weights[67][195] = 16'sd6;
        fc1_weights[67][196] = 16'sd-9;
        fc1_weights[67][197] = 16'sd-59;
        fc1_weights[67][198] = 16'sd-37;
        fc1_weights[67][199] = 16'sd-31;
        fc1_weights[67][200] = 16'sd-20;
        fc1_weights[67][201] = 16'sd-26;
        fc1_weights[67][202] = 16'sd-11;
        fc1_weights[67][203] = 16'sd-23;
        fc1_weights[67][204] = 16'sd-55;
        fc1_weights[67][205] = 16'sd-36;
        fc1_weights[67][206] = 16'sd13;
        fc1_weights[67][207] = 16'sd0;
        fc1_weights[68][0] = 16'sd105;
        fc1_weights[68][1] = 16'sd69;
        fc1_weights[68][2] = 16'sd71;
        fc1_weights[68][3] = 16'sd132;
        fc1_weights[68][4] = 16'sd83;
        fc1_weights[68][5] = 16'sd-10;
        fc1_weights[68][6] = 16'sd0;
        fc1_weights[68][7] = 16'sd39;
        fc1_weights[68][8] = 16'sd-61;
        fc1_weights[68][9] = 16'sd28;
        fc1_weights[68][10] = 16'sd-7;
        fc1_weights[68][11] = 16'sd30;
        fc1_weights[68][12] = 16'sd-29;
        fc1_weights[68][13] = 16'sd23;
        fc1_weights[68][14] = 16'sd84;
        fc1_weights[68][15] = 16'sd-7;
        fc1_weights[68][16] = 16'sd32;
        fc1_weights[68][17] = 16'sd-8;
        fc1_weights[68][18] = 16'sd35;
        fc1_weights[68][19] = 16'sd-41;
        fc1_weights[68][20] = 16'sd28;
        fc1_weights[68][21] = 16'sd23;
        fc1_weights[68][22] = 16'sd-13;
        fc1_weights[68][23] = 16'sd-39;
        fc1_weights[68][24] = 16'sd1;
        fc1_weights[68][25] = 16'sd-18;
        fc1_weights[68][26] = 16'sd19;
        fc1_weights[68][27] = 16'sd15;
        fc1_weights[68][28] = 16'sd56;
        fc1_weights[68][29] = 16'sd17;
        fc1_weights[68][30] = 16'sd-33;
        fc1_weights[68][31] = 16'sd-66;
        fc1_weights[68][32] = 16'sd-2;
        fc1_weights[68][33] = 16'sd103;
        fc1_weights[68][34] = 16'sd-4;
        fc1_weights[68][35] = 16'sd12;
        fc1_weights[68][36] = 16'sd63;
        fc1_weights[68][37] = 16'sd12;
        fc1_weights[68][38] = 16'sd-61;
        fc1_weights[68][39] = 16'sd68;
        fc1_weights[68][40] = 16'sd-12;
        fc1_weights[68][41] = 16'sd18;
        fc1_weights[68][42] = 16'sd48;
        fc1_weights[68][43] = 16'sd142;
        fc1_weights[68][44] = 16'sd56;
        fc1_weights[68][45] = 16'sd56;
        fc1_weights[68][46] = 16'sd98;
        fc1_weights[68][47] = 16'sd76;
        fc1_weights[68][48] = 16'sd36;
        fc1_weights[68][49] = 16'sd-28;
        fc1_weights[68][50] = 16'sd9;
        fc1_weights[68][51] = 16'sd-7;
        fc1_weights[68][52] = 16'sd-20;
        fc1_weights[68][53] = 16'sd40;
        fc1_weights[68][54] = 16'sd24;
        fc1_weights[68][55] = 16'sd7;
        fc1_weights[68][56] = 16'sd-61;
        fc1_weights[68][57] = 16'sd-47;
        fc1_weights[68][58] = 16'sd57;
        fc1_weights[68][59] = 16'sd23;
        fc1_weights[68][60] = 16'sd-84;
        fc1_weights[68][61] = 16'sd36;
        fc1_weights[68][62] = 16'sd38;
        fc1_weights[68][63] = 16'sd-19;
        fc1_weights[68][64] = 16'sd-49;
        fc1_weights[68][65] = 16'sd58;
        fc1_weights[68][66] = 16'sd-57;
        fc1_weights[68][67] = 16'sd2;
        fc1_weights[68][68] = 16'sd-27;
        fc1_weights[68][69] = 16'sd-61;
        fc1_weights[68][70] = 16'sd4;
        fc1_weights[68][71] = 16'sd-56;
        fc1_weights[68][72] = 16'sd-18;
        fc1_weights[68][73] = 16'sd-71;
        fc1_weights[68][74] = 16'sd-50;
        fc1_weights[68][75] = 16'sd-46;
        fc1_weights[68][76] = 16'sd-54;
        fc1_weights[68][77] = 16'sd-22;
        fc1_weights[68][78] = 16'sd-56;
        fc1_weights[68][79] = 16'sd10;
        fc1_weights[68][80] = 16'sd-12;
        fc1_weights[68][81] = 16'sd58;
        fc1_weights[68][82] = 16'sd79;
        fc1_weights[68][83] = 16'sd31;
        fc1_weights[68][84] = 16'sd90;
        fc1_weights[68][85] = 16'sd88;
        fc1_weights[68][86] = 16'sd11;
        fc1_weights[68][87] = 16'sd-42;
        fc1_weights[68][88] = 16'sd9;
        fc1_weights[68][89] = 16'sd-43;
        fc1_weights[68][90] = 16'sd-48;
        fc1_weights[68][91] = 16'sd-78;
        fc1_weights[68][92] = 16'sd-66;
        fc1_weights[68][93] = 16'sd34;
        fc1_weights[68][94] = 16'sd-12;
        fc1_weights[68][95] = 16'sd-66;
        fc1_weights[68][96] = 16'sd11;
        fc1_weights[68][97] = 16'sd-31;
        fc1_weights[68][98] = 16'sd-11;
        fc1_weights[68][99] = 16'sd-4;
        fc1_weights[68][100] = 16'sd-57;
        fc1_weights[68][101] = 16'sd24;
        fc1_weights[68][102] = 16'sd49;
        fc1_weights[68][103] = 16'sd-6;
        fc1_weights[68][104] = 16'sd-32;
        fc1_weights[68][105] = 16'sd2;
        fc1_weights[68][106] = 16'sd-2;
        fc1_weights[68][107] = 16'sd32;
        fc1_weights[68][108] = 16'sd-15;
        fc1_weights[68][109] = 16'sd-5;
        fc1_weights[68][110] = 16'sd-22;
        fc1_weights[68][111] = 16'sd-41;
        fc1_weights[68][112] = 16'sd-19;
        fc1_weights[68][113] = 16'sd11;
        fc1_weights[68][114] = 16'sd72;
        fc1_weights[68][115] = 16'sd24;
        fc1_weights[68][116] = 16'sd36;
        fc1_weights[68][117] = 16'sd-90;
        fc1_weights[68][118] = 16'sd-63;
        fc1_weights[68][119] = 16'sd-53;
        fc1_weights[68][120] = 16'sd-106;
        fc1_weights[68][121] = 16'sd-53;
        fc1_weights[68][122] = 16'sd27;
        fc1_weights[68][123] = 16'sd-45;
        fc1_weights[68][124] = 16'sd-15;
        fc1_weights[68][125] = 16'sd-8;
        fc1_weights[68][126] = 16'sd50;
        fc1_weights[68][127] = 16'sd2;
        fc1_weights[68][128] = 16'sd-22;
        fc1_weights[68][129] = 16'sd-14;
        fc1_weights[68][130] = 16'sd-37;
        fc1_weights[68][131] = 16'sd-52;
        fc1_weights[68][132] = 16'sd-96;
        fc1_weights[68][133] = 16'sd-75;
        fc1_weights[68][134] = 16'sd-15;
        fc1_weights[68][135] = 16'sd-50;
        fc1_weights[68][136] = 16'sd-67;
        fc1_weights[68][137] = 16'sd-9;
        fc1_weights[68][138] = 16'sd-8;
        fc1_weights[68][139] = 16'sd96;
        fc1_weights[68][140] = 16'sd48;
        fc1_weights[68][141] = 16'sd-17;
        fc1_weights[68][142] = 16'sd-94;
        fc1_weights[68][143] = 16'sd1;
        fc1_weights[68][144] = 16'sd-66;
        fc1_weights[68][145] = 16'sd38;
        fc1_weights[68][146] = 16'sd-15;
        fc1_weights[68][147] = 16'sd-65;
        fc1_weights[68][148] = 16'sd-25;
        fc1_weights[68][149] = 16'sd24;
        fc1_weights[68][150] = 16'sd-13;
        fc1_weights[68][151] = 16'sd32;
        fc1_weights[68][152] = 16'sd57;
        fc1_weights[68][153] = 16'sd39;
        fc1_weights[68][154] = 16'sd17;
        fc1_weights[68][155] = 16'sd33;
        fc1_weights[68][156] = 16'sd-11;
        fc1_weights[68][157] = 16'sd26;
        fc1_weights[68][158] = 16'sd-3;
        fc1_weights[68][159] = 16'sd46;
        fc1_weights[68][160] = 16'sd20;
        fc1_weights[68][161] = 16'sd-61;
        fc1_weights[68][162] = 16'sd-104;
        fc1_weights[68][163] = 16'sd-11;
        fc1_weights[68][164] = 16'sd36;
        fc1_weights[68][165] = 16'sd-15;
        fc1_weights[68][166] = 16'sd-27;
        fc1_weights[68][167] = 16'sd6;
        fc1_weights[68][168] = 16'sd-39;
        fc1_weights[68][169] = 16'sd-31;
        fc1_weights[68][170] = 16'sd-59;
        fc1_weights[68][171] = 16'sd-47;
        fc1_weights[68][172] = 16'sd33;
        fc1_weights[68][173] = 16'sd12;
        fc1_weights[68][174] = 16'sd-49;
        fc1_weights[68][175] = 16'sd4;
        fc1_weights[68][176] = 16'sd-18;
        fc1_weights[68][177] = 16'sd-22;
        fc1_weights[68][178] = 16'sd14;
        fc1_weights[68][179] = 16'sd34;
        fc1_weights[68][180] = 16'sd27;
        fc1_weights[68][181] = 16'sd70;
        fc1_weights[68][182] = 16'sd78;
        fc1_weights[68][183] = 16'sd28;
        fc1_weights[68][184] = 16'sd8;
        fc1_weights[68][185] = 16'sd-14;
        fc1_weights[68][186] = 16'sd45;
        fc1_weights[68][187] = 16'sd-21;
        fc1_weights[68][188] = 16'sd66;
        fc1_weights[68][189] = 16'sd18;
        fc1_weights[68][190] = 16'sd-27;
        fc1_weights[68][191] = 16'sd-24;
        fc1_weights[68][192] = 16'sd5;
        fc1_weights[68][193] = 16'sd4;
        fc1_weights[68][194] = 16'sd-58;
        fc1_weights[68][195] = 16'sd-38;
        fc1_weights[68][196] = 16'sd-17;
        fc1_weights[68][197] = 16'sd-37;
        fc1_weights[68][198] = 16'sd40;
        fc1_weights[68][199] = 16'sd40;
        fc1_weights[68][200] = 16'sd77;
        fc1_weights[68][201] = 16'sd51;
        fc1_weights[68][202] = 16'sd-40;
        fc1_weights[68][203] = 16'sd-37;
        fc1_weights[68][204] = 16'sd1;
        fc1_weights[68][205] = 16'sd42;
        fc1_weights[68][206] = 16'sd26;
        fc1_weights[68][207] = 16'sd63;
        fc1_weights[69][0] = 16'sd-19;
        fc1_weights[69][1] = 16'sd-8;
        fc1_weights[69][2] = 16'sd-105;
        fc1_weights[69][3] = 16'sd-8;
        fc1_weights[69][4] = 16'sd-40;
        fc1_weights[69][5] = 16'sd29;
        fc1_weights[69][6] = 16'sd54;
        fc1_weights[69][7] = 16'sd84;
        fc1_weights[69][8] = 16'sd-19;
        fc1_weights[69][9] = 16'sd25;
        fc1_weights[69][10] = 16'sd37;
        fc1_weights[69][11] = 16'sd-61;
        fc1_weights[69][12] = 16'sd-112;
        fc1_weights[69][13] = 16'sd-120;
        fc1_weights[69][14] = 16'sd-18;
        fc1_weights[69][15] = 16'sd40;
        fc1_weights[69][16] = 16'sd10;
        fc1_weights[69][17] = 16'sd-73;
        fc1_weights[69][18] = 16'sd-77;
        fc1_weights[69][19] = 16'sd-69;
        fc1_weights[69][20] = 16'sd28;
        fc1_weights[69][21] = 16'sd-29;
        fc1_weights[69][22] = 16'sd-6;
        fc1_weights[69][23] = 16'sd-47;
        fc1_weights[69][24] = 16'sd13;
        fc1_weights[69][25] = 16'sd-51;
        fc1_weights[69][26] = 16'sd-53;
        fc1_weights[69][27] = 16'sd-58;
        fc1_weights[69][28] = 16'sd-30;
        fc1_weights[69][29] = 16'sd-74;
        fc1_weights[69][30] = 16'sd4;
        fc1_weights[69][31] = 16'sd43;
        fc1_weights[69][32] = 16'sd-15;
        fc1_weights[69][33] = 16'sd17;
        fc1_weights[69][34] = 16'sd3;
        fc1_weights[69][35] = 16'sd8;
        fc1_weights[69][36] = 16'sd48;
        fc1_weights[69][37] = 16'sd37;
        fc1_weights[69][38] = 16'sd-48;
        fc1_weights[69][39] = 16'sd-109;
        fc1_weights[69][40] = 16'sd59;
        fc1_weights[69][41] = 16'sd44;
        fc1_weights[69][42] = 16'sd-17;
        fc1_weights[69][43] = 16'sd-10;
        fc1_weights[69][44] = 16'sd-33;
        fc1_weights[69][45] = 16'sd-108;
        fc1_weights[69][46] = 16'sd-25;
        fc1_weights[69][47] = 16'sd-5;
        fc1_weights[69][48] = 16'sd8;
        fc1_weights[69][49] = 16'sd-41;
        fc1_weights[69][50] = 16'sd-4;
        fc1_weights[69][51] = 16'sd-59;
        fc1_weights[69][52] = 16'sd-45;
        fc1_weights[69][53] = 16'sd-35;
        fc1_weights[69][54] = 16'sd29;
        fc1_weights[69][55] = 16'sd-50;
        fc1_weights[69][56] = 16'sd-53;
        fc1_weights[69][57] = 16'sd-3;
        fc1_weights[69][58] = 16'sd-31;
        fc1_weights[69][59] = 16'sd-16;
        fc1_weights[69][60] = 16'sd-18;
        fc1_weights[69][61] = 16'sd-7;
        fc1_weights[69][62] = 16'sd14;
        fc1_weights[69][63] = 16'sd9;
        fc1_weights[69][64] = 16'sd-39;
        fc1_weights[69][65] = 16'sd-23;
        fc1_weights[69][66] = 16'sd-27;
        fc1_weights[69][67] = 16'sd-6;
        fc1_weights[69][68] = 16'sd-62;
        fc1_weights[69][69] = 16'sd-105;
        fc1_weights[69][70] = 16'sd-69;
        fc1_weights[69][71] = 16'sd-14;
        fc1_weights[69][72] = 16'sd55;
        fc1_weights[69][73] = 16'sd-38;
        fc1_weights[69][74] = 16'sd25;
        fc1_weights[69][75] = 16'sd-20;
        fc1_weights[69][76] = 16'sd-6;
        fc1_weights[69][77] = 16'sd-72;
        fc1_weights[69][78] = 16'sd15;
        fc1_weights[69][79] = 16'sd67;
        fc1_weights[69][80] = 16'sd25;
        fc1_weights[69][81] = 16'sd42;
        fc1_weights[69][82] = 16'sd68;
        fc1_weights[69][83] = 16'sd62;
        fc1_weights[69][84] = 16'sd-6;
        fc1_weights[69][85] = 16'sd-50;
        fc1_weights[69][86] = 16'sd-58;
        fc1_weights[69][87] = 16'sd-39;
        fc1_weights[69][88] = 16'sd-79;
        fc1_weights[69][89] = 16'sd36;
        fc1_weights[69][90] = 16'sd-35;
        fc1_weights[69][91] = 16'sd-11;
        fc1_weights[69][92] = 16'sd46;
        fc1_weights[69][93] = 16'sd107;
        fc1_weights[69][94] = 16'sd2;
        fc1_weights[69][95] = 16'sd35;
        fc1_weights[69][96] = 16'sd-14;
        fc1_weights[69][97] = 16'sd-49;
        fc1_weights[69][98] = 16'sd2;
        fc1_weights[69][99] = 16'sd-10;
        fc1_weights[69][100] = 16'sd6;
        fc1_weights[69][101] = 16'sd9;
        fc1_weights[69][102] = 16'sd-3;
        fc1_weights[69][103] = 16'sd-47;
        fc1_weights[69][104] = 16'sd51;
        fc1_weights[69][105] = 16'sd-24;
        fc1_weights[69][106] = 16'sd12;
        fc1_weights[69][107] = 16'sd32;
        fc1_weights[69][108] = 16'sd-21;
        fc1_weights[69][109] = 16'sd-21;
        fc1_weights[69][110] = 16'sd-14;
        fc1_weights[69][111] = 16'sd-15;
        fc1_weights[69][112] = 16'sd6;
        fc1_weights[69][113] = 16'sd28;
        fc1_weights[69][114] = 16'sd-59;
        fc1_weights[69][115] = 16'sd-27;
        fc1_weights[69][116] = 16'sd42;
        fc1_weights[69][117] = 16'sd54;
        fc1_weights[69][118] = 16'sd42;
        fc1_weights[69][119] = 16'sd56;
        fc1_weights[69][120] = 16'sd21;
        fc1_weights[69][121] = 16'sd35;
        fc1_weights[69][122] = 16'sd52;
        fc1_weights[69][123] = 16'sd-9;
        fc1_weights[69][124] = 16'sd-47;
        fc1_weights[69][125] = 16'sd-36;
        fc1_weights[69][126] = 16'sd-62;
        fc1_weights[69][127] = 16'sd-7;
        fc1_weights[69][128] = 16'sd-42;
        fc1_weights[69][129] = 16'sd-117;
        fc1_weights[69][130] = 16'sd-27;
        fc1_weights[69][131] = 16'sd-43;
        fc1_weights[69][132] = 16'sd23;
        fc1_weights[69][133] = 16'sd-36;
        fc1_weights[69][134] = 16'sd-15;
        fc1_weights[69][135] = 16'sd20;
        fc1_weights[69][136] = 16'sd-4;
        fc1_weights[69][137] = 16'sd32;
        fc1_weights[69][138] = 16'sd-3;
        fc1_weights[69][139] = 16'sd22;
        fc1_weights[69][140] = 16'sd73;
        fc1_weights[69][141] = 16'sd-33;
        fc1_weights[69][142] = 16'sd107;
        fc1_weights[69][143] = 16'sd65;
        fc1_weights[69][144] = 16'sd62;
        fc1_weights[69][145] = 16'sd14;
        fc1_weights[69][146] = 16'sd11;
        fc1_weights[69][147] = 16'sd66;
        fc1_weights[69][148] = 16'sd45;
        fc1_weights[69][149] = 16'sd23;
        fc1_weights[69][150] = 16'sd5;
        fc1_weights[69][151] = 16'sd-9;
        fc1_weights[69][152] = 16'sd33;
        fc1_weights[69][153] = 16'sd22;
        fc1_weights[69][154] = 16'sd3;
        fc1_weights[69][155] = 16'sd28;
        fc1_weights[69][156] = 16'sd6;
        fc1_weights[69][157] = 16'sd29;
        fc1_weights[69][158] = 16'sd9;
        fc1_weights[69][159] = 16'sd25;
        fc1_weights[69][160] = 16'sd-15;
        fc1_weights[69][161] = 16'sd-42;
        fc1_weights[69][162] = 16'sd16;
        fc1_weights[69][163] = 16'sd-15;
        fc1_weights[69][164] = 16'sd26;
        fc1_weights[69][165] = 16'sd49;
        fc1_weights[69][166] = 16'sd101;
        fc1_weights[69][167] = 16'sd69;
        fc1_weights[69][168] = 16'sd44;
        fc1_weights[69][169] = 16'sd-30;
        fc1_weights[69][170] = 16'sd54;
        fc1_weights[69][171] = 16'sd22;
        fc1_weights[69][172] = 16'sd-8;
        fc1_weights[69][173] = 16'sd19;
        fc1_weights[69][174] = 16'sd-16;
        fc1_weights[69][175] = 16'sd6;
        fc1_weights[69][176] = 16'sd5;
        fc1_weights[69][177] = 16'sd18;
        fc1_weights[69][178] = 16'sd-22;
        fc1_weights[69][179] = 16'sd26;
        fc1_weights[69][180] = 16'sd22;
        fc1_weights[69][181] = 16'sd10;
        fc1_weights[69][182] = 16'sd-21;
        fc1_weights[69][183] = 16'sd10;
        fc1_weights[69][184] = 16'sd-24;
        fc1_weights[69][185] = 16'sd80;
        fc1_weights[69][186] = 16'sd-12;
        fc1_weights[69][187] = 16'sd-1;
        fc1_weights[69][188] = 16'sd11;
        fc1_weights[69][189] = 16'sd-4;
        fc1_weights[69][190] = 16'sd64;
        fc1_weights[69][191] = 16'sd101;
        fc1_weights[69][192] = 16'sd-17;
        fc1_weights[69][193] = 16'sd20;
        fc1_weights[69][194] = 16'sd27;
        fc1_weights[69][195] = 16'sd-5;
        fc1_weights[69][196] = 16'sd-8;
        fc1_weights[69][197] = 16'sd48;
        fc1_weights[69][198] = 16'sd1;
        fc1_weights[69][199] = 16'sd85;
        fc1_weights[69][200] = 16'sd-7;
        fc1_weights[69][201] = 16'sd19;
        fc1_weights[69][202] = 16'sd35;
        fc1_weights[69][203] = 16'sd-46;
        fc1_weights[69][204] = 16'sd-3;
        fc1_weights[69][205] = 16'sd31;
        fc1_weights[69][206] = 16'sd7;
        fc1_weights[69][207] = 16'sd-50;
        fc1_weights[70][0] = 16'sd32;
        fc1_weights[70][1] = 16'sd22;
        fc1_weights[70][2] = 16'sd85;
        fc1_weights[70][3] = 16'sd-24;
        fc1_weights[70][4] = 16'sd19;
        fc1_weights[70][5] = 16'sd36;
        fc1_weights[70][6] = 16'sd-2;
        fc1_weights[70][7] = 16'sd-38;
        fc1_weights[70][8] = 16'sd-48;
        fc1_weights[70][9] = 16'sd-80;
        fc1_weights[70][10] = 16'sd15;
        fc1_weights[70][11] = 16'sd5;
        fc1_weights[70][12] = 16'sd-27;
        fc1_weights[70][13] = 16'sd-19;
        fc1_weights[70][14] = 16'sd46;
        fc1_weights[70][15] = 16'sd15;
        fc1_weights[70][16] = 16'sd41;
        fc1_weights[70][17] = 16'sd49;
        fc1_weights[70][18] = 16'sd48;
        fc1_weights[70][19] = 16'sd11;
        fc1_weights[70][20] = 16'sd-44;
        fc1_weights[70][21] = 16'sd-28;
        fc1_weights[70][22] = 16'sd-63;
        fc1_weights[70][23] = 16'sd-16;
        fc1_weights[70][24] = 16'sd-36;
        fc1_weights[70][25] = 16'sd-37;
        fc1_weights[70][26] = 16'sd71;
        fc1_weights[70][27] = 16'sd54;
        fc1_weights[70][28] = 16'sd24;
        fc1_weights[70][29] = 16'sd20;
        fc1_weights[70][30] = 16'sd45;
        fc1_weights[70][31] = 16'sd72;
        fc1_weights[70][32] = 16'sd-7;
        fc1_weights[70][33] = 16'sd-50;
        fc1_weights[70][34] = 16'sd17;
        fc1_weights[70][35] = 16'sd-10;
        fc1_weights[70][36] = 16'sd-79;
        fc1_weights[70][37] = 16'sd27;
        fc1_weights[70][38] = 16'sd0;
        fc1_weights[70][39] = 16'sd34;
        fc1_weights[70][40] = 16'sd-34;
        fc1_weights[70][41] = 16'sd-13;
        fc1_weights[70][42] = 16'sd7;
        fc1_weights[70][43] = 16'sd11;
        fc1_weights[70][44] = 16'sd11;
        fc1_weights[70][45] = 16'sd-9;
        fc1_weights[70][46] = 16'sd-19;
        fc1_weights[70][47] = 16'sd-77;
        fc1_weights[70][48] = 16'sd-19;
        fc1_weights[70][49] = 16'sd-26;
        fc1_weights[70][50] = 16'sd24;
        fc1_weights[70][51] = 16'sd47;
        fc1_weights[70][52] = 16'sd12;
        fc1_weights[70][53] = 16'sd79;
        fc1_weights[70][54] = 16'sd7;
        fc1_weights[70][55] = 16'sd84;
        fc1_weights[70][56] = 16'sd89;
        fc1_weights[70][57] = 16'sd38;
        fc1_weights[70][58] = 16'sd31;
        fc1_weights[70][59] = 16'sd49;
        fc1_weights[70][60] = 16'sd-29;
        fc1_weights[70][61] = 16'sd-46;
        fc1_weights[70][62] = 16'sd-24;
        fc1_weights[70][63] = 16'sd-18;
        fc1_weights[70][64] = 16'sd-40;
        fc1_weights[70][65] = 16'sd-33;
        fc1_weights[70][66] = 16'sd-70;
        fc1_weights[70][67] = 16'sd3;
        fc1_weights[70][68] = 16'sd28;
        fc1_weights[70][69] = 16'sd-12;
        fc1_weights[70][70] = 16'sd43;
        fc1_weights[70][71] = 16'sd-55;
        fc1_weights[70][72] = 16'sd-43;
        fc1_weights[70][73] = 16'sd-34;
        fc1_weights[70][74] = 16'sd-77;
        fc1_weights[70][75] = 16'sd-16;
        fc1_weights[70][76] = 16'sd-6;
        fc1_weights[70][77] = 16'sd13;
        fc1_weights[70][78] = 16'sd-40;
        fc1_weights[70][79] = 16'sd-59;
        fc1_weights[70][80] = 16'sd89;
        fc1_weights[70][81] = 16'sd55;
        fc1_weights[70][82] = 16'sd20;
        fc1_weights[70][83] = 16'sd27;
        fc1_weights[70][84] = 16'sd-17;
        fc1_weights[70][85] = 16'sd7;
        fc1_weights[70][86] = 16'sd40;
        fc1_weights[70][87] = 16'sd44;
        fc1_weights[70][88] = 16'sd62;
        fc1_weights[70][89] = 16'sd-41;
        fc1_weights[70][90] = 16'sd-6;
        fc1_weights[70][91] = 16'sd-96;
        fc1_weights[70][92] = 16'sd-78;
        fc1_weights[70][93] = 16'sd-24;
        fc1_weights[70][94] = 16'sd3;
        fc1_weights[70][95] = 16'sd9;
        fc1_weights[70][96] = 16'sd-2;
        fc1_weights[70][97] = 16'sd18;
        fc1_weights[70][98] = 16'sd-49;
        fc1_weights[70][99] = 16'sd6;
        fc1_weights[70][100] = 16'sd-91;
        fc1_weights[70][101] = 16'sd-39;
        fc1_weights[70][102] = 16'sd-32;
        fc1_weights[70][103] = 16'sd1;
        fc1_weights[70][104] = 16'sd7;
        fc1_weights[70][105] = 16'sd-7;
        fc1_weights[70][106] = 16'sd6;
        fc1_weights[70][107] = 16'sd3;
        fc1_weights[70][108] = 16'sd17;
        fc1_weights[70][109] = 16'sd33;
        fc1_weights[70][110] = 16'sd6;
        fc1_weights[70][111] = 16'sd36;
        fc1_weights[70][112] = 16'sd11;
        fc1_weights[70][113] = 16'sd45;
        fc1_weights[70][114] = 16'sd-50;
        fc1_weights[70][115] = 16'sd13;
        fc1_weights[70][116] = 16'sd-111;
        fc1_weights[70][117] = 16'sd-40;
        fc1_weights[70][118] = 16'sd23;
        fc1_weights[70][119] = 16'sd-35;
        fc1_weights[70][120] = 16'sd-32;
        fc1_weights[70][121] = 16'sd-38;
        fc1_weights[70][122] = 16'sd-72;
        fc1_weights[70][123] = 16'sd-50;
        fc1_weights[70][124] = 16'sd-32;
        fc1_weights[70][125] = 16'sd-42;
        fc1_weights[70][126] = 16'sd-19;
        fc1_weights[70][127] = 16'sd14;
        fc1_weights[70][128] = 16'sd16;
        fc1_weights[70][129] = 16'sd25;
        fc1_weights[70][130] = 16'sd-7;
        fc1_weights[70][131] = 16'sd-31;
        fc1_weights[70][132] = 16'sd-10;
        fc1_weights[70][133] = 16'sd58;
        fc1_weights[70][134] = 16'sd-31;
        fc1_weights[70][135] = 16'sd-7;
        fc1_weights[70][136] = 16'sd28;
        fc1_weights[70][137] = 16'sd-14;
        fc1_weights[70][138] = 16'sd55;
        fc1_weights[70][139] = 16'sd-33;
        fc1_weights[70][140] = 16'sd-84;
        fc1_weights[70][141] = 16'sd11;
        fc1_weights[70][142] = 16'sd-73;
        fc1_weights[70][143] = 16'sd15;
        fc1_weights[70][144] = 16'sd24;
        fc1_weights[70][145] = 16'sd51;
        fc1_weights[70][146] = 16'sd7;
        fc1_weights[70][147] = 16'sd-8;
        fc1_weights[70][148] = 16'sd-5;
        fc1_weights[70][149] = 16'sd-48;
        fc1_weights[70][150] = 16'sd-38;
        fc1_weights[70][151] = 16'sd-20;
        fc1_weights[70][152] = 16'sd-18;
        fc1_weights[70][153] = 16'sd-29;
        fc1_weights[70][154] = 16'sd-81;
        fc1_weights[70][155] = 16'sd-6;
        fc1_weights[70][156] = 16'sd-37;
        fc1_weights[70][157] = 16'sd-10;
        fc1_weights[70][158] = 16'sd7;
        fc1_weights[70][159] = 16'sd-30;
        fc1_weights[70][160] = 16'sd-5;
        fc1_weights[70][161] = 16'sd45;
        fc1_weights[70][162] = 16'sd53;
        fc1_weights[70][163] = 16'sd18;
        fc1_weights[70][164] = 16'sd-5;
        fc1_weights[70][165] = 16'sd-8;
        fc1_weights[70][166] = 16'sd-62;
        fc1_weights[70][167] = 16'sd-72;
        fc1_weights[70][168] = 16'sd-46;
        fc1_weights[70][169] = 16'sd7;
        fc1_weights[70][170] = 16'sd49;
        fc1_weights[70][171] = 16'sd-39;
        fc1_weights[70][172] = 16'sd16;
        fc1_weights[70][173] = 16'sd-35;
        fc1_weights[70][174] = 16'sd-13;
        fc1_weights[70][175] = 16'sd-33;
        fc1_weights[70][176] = 16'sd16;
        fc1_weights[70][177] = 16'sd34;
        fc1_weights[70][178] = 16'sd-21;
        fc1_weights[70][179] = 16'sd-47;
        fc1_weights[70][180] = 16'sd-18;
        fc1_weights[70][181] = 16'sd-28;
        fc1_weights[70][182] = 16'sd-25;
        fc1_weights[70][183] = 16'sd-60;
        fc1_weights[70][184] = 16'sd14;
        fc1_weights[70][185] = 16'sd-7;
        fc1_weights[70][186] = 16'sd95;
        fc1_weights[70][187] = 16'sd11;
        fc1_weights[70][188] = 16'sd25;
        fc1_weights[70][189] = 16'sd69;
        fc1_weights[70][190] = 16'sd85;
        fc1_weights[70][191] = 16'sd-19;
        fc1_weights[70][192] = 16'sd57;
        fc1_weights[70][193] = 16'sd27;
        fc1_weights[70][194] = 16'sd52;
        fc1_weights[70][195] = 16'sd35;
        fc1_weights[70][196] = 16'sd92;
        fc1_weights[70][197] = 16'sd36;
        fc1_weights[70][198] = 16'sd46;
        fc1_weights[70][199] = 16'sd70;
        fc1_weights[70][200] = 16'sd24;
        fc1_weights[70][201] = 16'sd20;
        fc1_weights[70][202] = 16'sd3;
        fc1_weights[70][203] = 16'sd31;
        fc1_weights[70][204] = 16'sd8;
        fc1_weights[70][205] = 16'sd-42;
        fc1_weights[70][206] = 16'sd41;
        fc1_weights[70][207] = 16'sd43;
        fc1_weights[71][0] = 16'sd-21;
        fc1_weights[71][1] = 16'sd29;
        fc1_weights[71][2] = 16'sd17;
        fc1_weights[71][3] = 16'sd17;
        fc1_weights[71][4] = 16'sd-35;
        fc1_weights[71][5] = 16'sd-10;
        fc1_weights[71][6] = 16'sd-11;
        fc1_weights[71][7] = 16'sd-71;
        fc1_weights[71][8] = 16'sd-34;
        fc1_weights[71][9] = 16'sd39;
        fc1_weights[71][10] = 16'sd10;
        fc1_weights[71][11] = 16'sd15;
        fc1_weights[71][12] = 16'sd3;
        fc1_weights[71][13] = 16'sd44;
        fc1_weights[71][14] = 16'sd-10;
        fc1_weights[71][15] = 16'sd40;
        fc1_weights[71][16] = 16'sd14;
        fc1_weights[71][17] = 16'sd-43;
        fc1_weights[71][18] = 16'sd-22;
        fc1_weights[71][19] = 16'sd-51;
        fc1_weights[71][20] = 16'sd9;
        fc1_weights[71][21] = 16'sd14;
        fc1_weights[71][22] = 16'sd30;
        fc1_weights[71][23] = 16'sd18;
        fc1_weights[71][24] = 16'sd64;
        fc1_weights[71][25] = 16'sd67;
        fc1_weights[71][26] = 16'sd-5;
        fc1_weights[71][27] = 16'sd7;
        fc1_weights[71][28] = 16'sd-13;
        fc1_weights[71][29] = 16'sd21;
        fc1_weights[71][30] = 16'sd-2;
        fc1_weights[71][31] = 16'sd-46;
        fc1_weights[71][32] = 16'sd-10;
        fc1_weights[71][33] = 16'sd-106;
        fc1_weights[71][34] = 16'sd-7;
        fc1_weights[71][35] = 16'sd-46;
        fc1_weights[71][36] = 16'sd33;
        fc1_weights[71][37] = 16'sd-59;
        fc1_weights[71][38] = 16'sd-8;
        fc1_weights[71][39] = 16'sd38;
        fc1_weights[71][40] = 16'sd97;
        fc1_weights[71][41] = 16'sd63;
        fc1_weights[71][42] = 16'sd-59;
        fc1_weights[71][43] = 16'sd2;
        fc1_weights[71][44] = 16'sd24;
        fc1_weights[71][45] = 16'sd-3;
        fc1_weights[71][46] = 16'sd20;
        fc1_weights[71][47] = 16'sd-3;
        fc1_weights[71][48] = 16'sd-64;
        fc1_weights[71][49] = 16'sd31;
        fc1_weights[71][50] = 16'sd30;
        fc1_weights[71][51] = 16'sd22;
        fc1_weights[71][52] = 16'sd20;
        fc1_weights[71][53] = 16'sd36;
        fc1_weights[71][54] = 16'sd-45;
        fc1_weights[71][55] = 16'sd-12;
        fc1_weights[71][56] = 16'sd20;
        fc1_weights[71][57] = 16'sd-47;
        fc1_weights[71][58] = 16'sd-31;
        fc1_weights[71][59] = 16'sd-45;
        fc1_weights[71][60] = 16'sd22;
        fc1_weights[71][61] = 16'sd-33;
        fc1_weights[71][62] = 16'sd-20;
        fc1_weights[71][63] = 16'sd13;
        fc1_weights[71][64] = 16'sd24;
        fc1_weights[71][65] = 16'sd30;
        fc1_weights[71][66] = 16'sd71;
        fc1_weights[71][67] = 16'sd-37;
        fc1_weights[71][68] = 16'sd-61;
        fc1_weights[71][69] = 16'sd-13;
        fc1_weights[71][70] = 16'sd48;
        fc1_weights[71][71] = 16'sd42;
        fc1_weights[71][72] = 16'sd-44;
        fc1_weights[71][73] = 16'sd-25;
        fc1_weights[71][74] = 16'sd10;
        fc1_weights[71][75] = 16'sd-11;
        fc1_weights[71][76] = 16'sd29;
        fc1_weights[71][77] = 16'sd45;
        fc1_weights[71][78] = 16'sd44;
        fc1_weights[71][79] = 16'sd76;
        fc1_weights[71][80] = 16'sd10;
        fc1_weights[71][81] = 16'sd-4;
        fc1_weights[71][82] = 16'sd-30;
        fc1_weights[71][83] = 16'sd-65;
        fc1_weights[71][84] = 16'sd-44;
        fc1_weights[71][85] = 16'sd-48;
        fc1_weights[71][86] = 16'sd3;
        fc1_weights[71][87] = 16'sd51;
        fc1_weights[71][88] = 16'sd61;
        fc1_weights[71][89] = 16'sd7;
        fc1_weights[71][90] = 16'sd122;
        fc1_weights[71][91] = 16'sd98;
        fc1_weights[71][92] = 16'sd59;
        fc1_weights[71][93] = 16'sd-9;
        fc1_weights[71][94] = 16'sd-45;
        fc1_weights[71][95] = 16'sd-24;
        fc1_weights[71][96] = 16'sd-10;
        fc1_weights[71][97] = 16'sd33;
        fc1_weights[71][98] = 16'sd-32;
        fc1_weights[71][99] = 16'sd-19;
        fc1_weights[71][100] = 16'sd-24;
        fc1_weights[71][101] = 16'sd0;
        fc1_weights[71][102] = 16'sd17;
        fc1_weights[71][103] = 16'sd29;
        fc1_weights[71][104] = 16'sd25;
        fc1_weights[71][105] = 16'sd18;
        fc1_weights[71][106] = 16'sd-2;
        fc1_weights[71][107] = 16'sd13;
        fc1_weights[71][108] = 16'sd-7;
        fc1_weights[71][109] = 16'sd-38;
        fc1_weights[71][110] = 16'sd-45;
        fc1_weights[71][111] = 16'sd14;
        fc1_weights[71][112] = 16'sd28;
        fc1_weights[71][113] = 16'sd-24;
        fc1_weights[71][114] = 16'sd4;
        fc1_weights[71][115] = 16'sd-32;
        fc1_weights[71][116] = 16'sd47;
        fc1_weights[71][117] = 16'sd18;
        fc1_weights[71][118] = 16'sd33;
        fc1_weights[71][119] = 16'sd20;
        fc1_weights[71][120] = 16'sd34;
        fc1_weights[71][121] = 16'sd49;
        fc1_weights[71][122] = 16'sd62;
        fc1_weights[71][123] = 16'sd43;
        fc1_weights[71][124] = 16'sd-32;
        fc1_weights[71][125] = 16'sd24;
        fc1_weights[71][126] = 16'sd-28;
        fc1_weights[71][127] = 16'sd-4;
        fc1_weights[71][128] = 16'sd-2;
        fc1_weights[71][129] = 16'sd-2;
        fc1_weights[71][130] = 16'sd-22;
        fc1_weights[71][131] = 16'sd19;
        fc1_weights[71][132] = 16'sd24;
        fc1_weights[71][133] = 16'sd38;
        fc1_weights[71][134] = 16'sd50;
        fc1_weights[71][135] = 16'sd48;
        fc1_weights[71][136] = 16'sd47;
        fc1_weights[71][137] = 16'sd12;
        fc1_weights[71][138] = 16'sd-19;
        fc1_weights[71][139] = 16'sd-63;
        fc1_weights[71][140] = 16'sd-78;
        fc1_weights[71][141] = 16'sd-99;
        fc1_weights[71][142] = 16'sd10;
        fc1_weights[71][143] = 16'sd4;
        fc1_weights[71][144] = 16'sd8;
        fc1_weights[71][145] = 16'sd-64;
        fc1_weights[71][146] = 16'sd-30;
        fc1_weights[71][147] = 16'sd6;
        fc1_weights[71][148] = 16'sd-14;
        fc1_weights[71][149] = 16'sd-26;
        fc1_weights[71][150] = 16'sd-1;
        fc1_weights[71][151] = 16'sd17;
        fc1_weights[71][152] = 16'sd-26;
        fc1_weights[71][153] = 16'sd-25;
        fc1_weights[71][154] = 16'sd-14;
        fc1_weights[71][155] = 16'sd22;
        fc1_weights[71][156] = 16'sd6;
        fc1_weights[71][157] = 16'sd20;
        fc1_weights[71][158] = 16'sd40;
        fc1_weights[71][159] = 16'sd-22;
        fc1_weights[71][160] = 16'sd-38;
        fc1_weights[71][161] = 16'sd-22;
        fc1_weights[71][162] = 16'sd21;
        fc1_weights[71][163] = 16'sd-14;
        fc1_weights[71][164] = 16'sd-57;
        fc1_weights[71][165] = 16'sd-39;
        fc1_weights[71][166] = 16'sd1;
        fc1_weights[71][167] = 16'sd8;
        fc1_weights[71][168] = 16'sd-8;
        fc1_weights[71][169] = 16'sd-17;
        fc1_weights[71][170] = 16'sd17;
        fc1_weights[71][171] = 16'sd-67;
        fc1_weights[71][172] = 16'sd-29;
        fc1_weights[71][173] = 16'sd-22;
        fc1_weights[71][174] = 16'sd-11;
        fc1_weights[71][175] = 16'sd-35;
        fc1_weights[71][176] = 16'sd-25;
        fc1_weights[71][177] = 16'sd-6;
        fc1_weights[71][178] = 16'sd-26;
        fc1_weights[71][179] = 16'sd16;
        fc1_weights[71][180] = 16'sd4;
        fc1_weights[71][181] = 16'sd36;
        fc1_weights[71][182] = 16'sd-17;
        fc1_weights[71][183] = 16'sd-18;
        fc1_weights[71][184] = 16'sd-15;
        fc1_weights[71][185] = 16'sd-42;
        fc1_weights[71][186] = 16'sd0;
        fc1_weights[71][187] = 16'sd20;
        fc1_weights[71][188] = 16'sd20;
        fc1_weights[71][189] = 16'sd-7;
        fc1_weights[71][190] = 16'sd-4;
        fc1_weights[71][191] = 16'sd41;
        fc1_weights[71][192] = 16'sd17;
        fc1_weights[71][193] = 16'sd1;
        fc1_weights[71][194] = 16'sd-9;
        fc1_weights[71][195] = 16'sd-4;
        fc1_weights[71][196] = 16'sd1;
        fc1_weights[71][197] = 16'sd82;
        fc1_weights[71][198] = 16'sd-24;
        fc1_weights[71][199] = 16'sd-47;
        fc1_weights[71][200] = 16'sd9;
        fc1_weights[71][201] = 16'sd-18;
        fc1_weights[71][202] = 16'sd-32;
        fc1_weights[71][203] = 16'sd48;
        fc1_weights[71][204] = 16'sd20;
        fc1_weights[71][205] = 16'sd-11;
        fc1_weights[71][206] = 16'sd-30;
        fc1_weights[71][207] = 16'sd-8;
        fc1_weights[72][0] = 16'sd19;
        fc1_weights[72][1] = 16'sd23;
        fc1_weights[72][2] = 16'sd70;
        fc1_weights[72][3] = 16'sd4;
        fc1_weights[72][4] = 16'sd58;
        fc1_weights[72][5] = 16'sd14;
        fc1_weights[72][6] = 16'sd43;
        fc1_weights[72][7] = 16'sd-31;
        fc1_weights[72][8] = 16'sd-16;
        fc1_weights[72][9] = 16'sd10;
        fc1_weights[72][10] = 16'sd20;
        fc1_weights[72][11] = 16'sd-7;
        fc1_weights[72][12] = 16'sd44;
        fc1_weights[72][13] = 16'sd66;
        fc1_weights[72][14] = 16'sd76;
        fc1_weights[72][15] = 16'sd37;
        fc1_weights[72][16] = 16'sd6;
        fc1_weights[72][17] = 16'sd44;
        fc1_weights[72][18] = 16'sd44;
        fc1_weights[72][19] = 16'sd59;
        fc1_weights[72][20] = 16'sd6;
        fc1_weights[72][21] = 16'sd3;
        fc1_weights[72][22] = 16'sd30;
        fc1_weights[72][23] = 16'sd94;
        fc1_weights[72][24] = 16'sd-14;
        fc1_weights[72][25] = 16'sd5;
        fc1_weights[72][26] = 16'sd63;
        fc1_weights[72][27] = 16'sd-24;
        fc1_weights[72][28] = 16'sd-3;
        fc1_weights[72][29] = 16'sd-38;
        fc1_weights[72][30] = 16'sd-18;
        fc1_weights[72][31] = 16'sd8;
        fc1_weights[72][32] = 16'sd16;
        fc1_weights[72][33] = 16'sd22;
        fc1_weights[72][34] = 16'sd-51;
        fc1_weights[72][35] = 16'sd-31;
        fc1_weights[72][36] = 16'sd-19;
        fc1_weights[72][37] = 16'sd1;
        fc1_weights[72][38] = 16'sd14;
        fc1_weights[72][39] = 16'sd41;
        fc1_weights[72][40] = 16'sd-28;
        fc1_weights[72][41] = 16'sd-64;
        fc1_weights[72][42] = 16'sd36;
        fc1_weights[72][43] = 16'sd59;
        fc1_weights[72][44] = 16'sd74;
        fc1_weights[72][45] = 16'sd21;
        fc1_weights[72][46] = 16'sd2;
        fc1_weights[72][47] = 16'sd31;
        fc1_weights[72][48] = 16'sd48;
        fc1_weights[72][49] = 16'sd-27;
        fc1_weights[72][50] = 16'sd12;
        fc1_weights[72][51] = 16'sd-28;
        fc1_weights[72][52] = 16'sd82;
        fc1_weights[72][53] = 16'sd-1;
        fc1_weights[72][54] = 16'sd13;
        fc1_weights[72][55] = 16'sd4;
        fc1_weights[72][56] = 16'sd0;
        fc1_weights[72][57] = 16'sd35;
        fc1_weights[72][58] = 16'sd-23;
        fc1_weights[72][59] = 16'sd1;
        fc1_weights[72][60] = 16'sd-20;
        fc1_weights[72][61] = 16'sd-10;
        fc1_weights[72][62] = 16'sd16;
        fc1_weights[72][63] = 16'sd-35;
        fc1_weights[72][64] = 16'sd-65;
        fc1_weights[72][65] = 16'sd-49;
        fc1_weights[72][66] = 16'sd-38;
        fc1_weights[72][67] = 16'sd-4;
        fc1_weights[72][68] = 16'sd57;
        fc1_weights[72][69] = 16'sd-8;
        fc1_weights[72][70] = 16'sd28;
        fc1_weights[72][71] = 16'sd-72;
        fc1_weights[72][72] = 16'sd-18;
        fc1_weights[72][73] = 16'sd15;
        fc1_weights[72][74] = 16'sd19;
        fc1_weights[72][75] = 16'sd-29;
        fc1_weights[72][76] = 16'sd-31;
        fc1_weights[72][77] = 16'sd-88;
        fc1_weights[72][78] = 16'sd55;
        fc1_weights[72][79] = 16'sd-29;
        fc1_weights[72][80] = 16'sd45;
        fc1_weights[72][81] = 16'sd37;
        fc1_weights[72][82] = 16'sd42;
        fc1_weights[72][83] = 16'sd13;
        fc1_weights[72][84] = 16'sd45;
        fc1_weights[72][85] = 16'sd76;
        fc1_weights[72][86] = 16'sd74;
        fc1_weights[72][87] = 16'sd40;
        fc1_weights[72][88] = 16'sd65;
        fc1_weights[72][89] = 16'sd-69;
        fc1_weights[72][90] = 16'sd-61;
        fc1_weights[72][91] = 16'sd22;
        fc1_weights[72][92] = 16'sd-10;
        fc1_weights[72][93] = 16'sd9;
        fc1_weights[72][94] = 16'sd51;
        fc1_weights[72][95] = 16'sd-61;
        fc1_weights[72][96] = 16'sd16;
        fc1_weights[72][97] = 16'sd-59;
        fc1_weights[72][98] = 16'sd-41;
        fc1_weights[72][99] = 16'sd33;
        fc1_weights[72][100] = 16'sd1;
        fc1_weights[72][101] = 16'sd5;
        fc1_weights[72][102] = 16'sd8;
        fc1_weights[72][103] = 16'sd2;
        fc1_weights[72][104] = 16'sd-23;
        fc1_weights[72][105] = 16'sd4;
        fc1_weights[72][106] = 16'sd9;
        fc1_weights[72][107] = 16'sd-8;
        fc1_weights[72][108] = 16'sd-7;
        fc1_weights[72][109] = 16'sd5;
        fc1_weights[72][110] = 16'sd57;
        fc1_weights[72][111] = 16'sd88;
        fc1_weights[72][112] = 16'sd-52;
        fc1_weights[72][113] = 16'sd-69;
        fc1_weights[72][114] = 16'sd2;
        fc1_weights[72][115] = 16'sd1;
        fc1_weights[72][116] = 16'sd22;
        fc1_weights[72][117] = 16'sd-43;
        fc1_weights[72][118] = 16'sd-42;
        fc1_weights[72][119] = 16'sd-28;
        fc1_weights[72][120] = 16'sd-32;
        fc1_weights[72][121] = 16'sd-25;
        fc1_weights[72][122] = 16'sd16;
        fc1_weights[72][123] = 16'sd37;
        fc1_weights[72][124] = 16'sd108;
        fc1_weights[72][125] = 16'sd99;
        fc1_weights[72][126] = 16'sd51;
        fc1_weights[72][127] = 16'sd22;
        fc1_weights[72][128] = 16'sd-5;
        fc1_weights[72][129] = 16'sd61;
        fc1_weights[72][130] = 16'sd-8;
        fc1_weights[72][131] = 16'sd32;
        fc1_weights[72][132] = 16'sd-14;
        fc1_weights[72][133] = 16'sd16;
        fc1_weights[72][134] = 16'sd-16;
        fc1_weights[72][135] = 16'sd-47;
        fc1_weights[72][136] = 16'sd61;
        fc1_weights[72][137] = 16'sd32;
        fc1_weights[72][138] = 16'sd42;
        fc1_weights[72][139] = 16'sd24;
        fc1_weights[72][140] = 16'sd26;
        fc1_weights[72][141] = 16'sd93;
        fc1_weights[72][142] = 16'sd-32;
        fc1_weights[72][143] = 16'sd82;
        fc1_weights[72][144] = 16'sd22;
        fc1_weights[72][145] = 16'sd62;
        fc1_weights[72][146] = 16'sd25;
        fc1_weights[72][147] = 16'sd19;
        fc1_weights[72][148] = 16'sd65;
        fc1_weights[72][149] = 16'sd14;
        fc1_weights[72][150] = 16'sd62;
        fc1_weights[72][151] = 16'sd28;
        fc1_weights[72][152] = 16'sd26;
        fc1_weights[72][153] = 16'sd-42;
        fc1_weights[72][154] = 16'sd-5;
        fc1_weights[72][155] = 16'sd14;
        fc1_weights[72][156] = 16'sd7;
        fc1_weights[72][157] = 16'sd15;
        fc1_weights[72][158] = 16'sd3;
        fc1_weights[72][159] = 16'sd-34;
        fc1_weights[72][160] = 16'sd17;
        fc1_weights[72][161] = 16'sd29;
        fc1_weights[72][162] = 16'sd1;
        fc1_weights[72][163] = 16'sd11;
        fc1_weights[72][164] = 16'sd60;
        fc1_weights[72][165] = 16'sd55;
        fc1_weights[72][166] = 16'sd44;
        fc1_weights[72][167] = 16'sd-4;
        fc1_weights[72][168] = 16'sd-32;
        fc1_weights[72][169] = 16'sd-19;
        fc1_weights[72][170] = 16'sd-68;
        fc1_weights[72][171] = 16'sd-75;
        fc1_weights[72][172] = 16'sd-28;
        fc1_weights[72][173] = 16'sd-36;
        fc1_weights[72][174] = 16'sd-5;
        fc1_weights[72][175] = 16'sd-18;
        fc1_weights[72][176] = 16'sd6;
        fc1_weights[72][177] = 16'sd15;
        fc1_weights[72][178] = 16'sd42;
        fc1_weights[72][179] = 16'sd10;
        fc1_weights[72][180] = 16'sd-2;
        fc1_weights[72][181] = 16'sd24;
        fc1_weights[72][182] = 16'sd-54;
        fc1_weights[72][183] = 16'sd-13;
        fc1_weights[72][184] = 16'sd-30;
        fc1_weights[72][185] = 16'sd-86;
        fc1_weights[72][186] = 16'sd-61;
        fc1_weights[72][187] = 16'sd-15;
        fc1_weights[72][188] = 16'sd-44;
        fc1_weights[72][189] = 16'sd14;
        fc1_weights[72][190] = 16'sd25;
        fc1_weights[72][191] = 16'sd9;
        fc1_weights[72][192] = 16'sd0;
        fc1_weights[72][193] = 16'sd28;
        fc1_weights[72][194] = 16'sd-3;
        fc1_weights[72][195] = 16'sd-18;
        fc1_weights[72][196] = 16'sd-11;
        fc1_weights[72][197] = 16'sd-39;
        fc1_weights[72][198] = 16'sd-80;
        fc1_weights[72][199] = 16'sd-33;
        fc1_weights[72][200] = 16'sd-44;
        fc1_weights[72][201] = 16'sd-30;
        fc1_weights[72][202] = 16'sd-8;
        fc1_weights[72][203] = 16'sd-1;
        fc1_weights[72][204] = 16'sd19;
        fc1_weights[72][205] = 16'sd1;
        fc1_weights[72][206] = 16'sd50;
        fc1_weights[72][207] = 16'sd3;
        fc1_weights[73][0] = 16'sd14;
        fc1_weights[73][1] = 16'sd25;
        fc1_weights[73][2] = 16'sd2;
        fc1_weights[73][3] = 16'sd68;
        fc1_weights[73][4] = 16'sd16;
        fc1_weights[73][5] = 16'sd5;
        fc1_weights[73][6] = 16'sd7;
        fc1_weights[73][7] = 16'sd28;
        fc1_weights[73][8] = 16'sd6;
        fc1_weights[73][9] = 16'sd-1;
        fc1_weights[73][10] = 16'sd-11;
        fc1_weights[73][11] = 16'sd66;
        fc1_weights[73][12] = 16'sd66;
        fc1_weights[73][13] = 16'sd-12;
        fc1_weights[73][14] = 16'sd-1;
        fc1_weights[73][15] = 16'sd15;
        fc1_weights[73][16] = 16'sd22;
        fc1_weights[73][17] = 16'sd32;
        fc1_weights[73][18] = 16'sd31;
        fc1_weights[73][19] = 16'sd47;
        fc1_weights[73][20] = 16'sd6;
        fc1_weights[73][21] = 16'sd-4;
        fc1_weights[73][22] = 16'sd-36;
        fc1_weights[73][23] = 16'sd-9;
        fc1_weights[73][24] = 16'sd-48;
        fc1_weights[73][25] = 16'sd-59;
        fc1_weights[73][26] = 16'sd-75;
        fc1_weights[73][27] = 16'sd-13;
        fc1_weights[73][28] = 16'sd-21;
        fc1_weights[73][29] = 16'sd19;
        fc1_weights[73][30] = 16'sd-41;
        fc1_weights[73][31] = 16'sd-15;
        fc1_weights[73][32] = 16'sd-17;
        fc1_weights[73][33] = 16'sd55;
        fc1_weights[73][34] = 16'sd29;
        fc1_weights[73][35] = 16'sd-24;
        fc1_weights[73][36] = 16'sd-32;
        fc1_weights[73][37] = 16'sd-4;
        fc1_weights[73][38] = 16'sd39;
        fc1_weights[73][39] = 16'sd28;
        fc1_weights[73][40] = 16'sd-12;
        fc1_weights[73][41] = 16'sd36;
        fc1_weights[73][42] = 16'sd92;
        fc1_weights[73][43] = 16'sd23;
        fc1_weights[73][44] = 16'sd16;
        fc1_weights[73][45] = 16'sd57;
        fc1_weights[73][46] = 16'sd-8;
        fc1_weights[73][47] = 16'sd-21;
        fc1_weights[73][48] = 16'sd-33;
        fc1_weights[73][49] = 16'sd-31;
        fc1_weights[73][50] = 16'sd-23;
        fc1_weights[73][51] = 16'sd-19;
        fc1_weights[73][52] = 16'sd-63;
        fc1_weights[73][53] = 16'sd-5;
        fc1_weights[73][54] = 16'sd23;
        fc1_weights[73][55] = 16'sd-40;
        fc1_weights[73][56] = 16'sd-63;
        fc1_weights[73][57] = 16'sd-42;
        fc1_weights[73][58] = 16'sd-33;
        fc1_weights[73][59] = 16'sd10;
        fc1_weights[73][60] = 16'sd65;
        fc1_weights[73][61] = 16'sd-3;
        fc1_weights[73][62] = 16'sd47;
        fc1_weights[73][63] = 16'sd-41;
        fc1_weights[73][64] = 16'sd30;
        fc1_weights[73][65] = 16'sd17;
        fc1_weights[73][66] = 16'sd10;
        fc1_weights[73][67] = 16'sd-4;
        fc1_weights[73][68] = 16'sd1;
        fc1_weights[73][69] = 16'sd68;
        fc1_weights[73][70] = 16'sd-14;
        fc1_weights[73][71] = 16'sd-4;
        fc1_weights[73][72] = 16'sd-2;
        fc1_weights[73][73] = 16'sd1;
        fc1_weights[73][74] = 16'sd-28;
        fc1_weights[73][75] = 16'sd-3;
        fc1_weights[73][76] = 16'sd-18;
        fc1_weights[73][77] = 16'sd23;
        fc1_weights[73][78] = 16'sd-36;
        fc1_weights[73][79] = 16'sd-92;
        fc1_weights[73][80] = 16'sd-64;
        fc1_weights[73][81] = 16'sd-40;
        fc1_weights[73][82] = 16'sd2;
        fc1_weights[73][83] = 16'sd21;
        fc1_weights[73][84] = 16'sd36;
        fc1_weights[73][85] = 16'sd41;
        fc1_weights[73][86] = 16'sd56;
        fc1_weights[73][87] = 16'sd-64;
        fc1_weights[73][88] = 16'sd-50;
        fc1_weights[73][89] = 16'sd37;
        fc1_weights[73][90] = 16'sd11;
        fc1_weights[73][91] = 16'sd-14;
        fc1_weights[73][92] = 16'sd-7;
        fc1_weights[73][93] = 16'sd-74;
        fc1_weights[73][94] = 16'sd50;
        fc1_weights[73][95] = 16'sd9;
        fc1_weights[73][96] = 16'sd28;
        fc1_weights[73][97] = 16'sd-7;
        fc1_weights[73][98] = 16'sd-24;
        fc1_weights[73][99] = 16'sd0;
        fc1_weights[73][100] = 16'sd-40;
        fc1_weights[73][101] = 16'sd42;
        fc1_weights[73][102] = 16'sd16;
        fc1_weights[73][103] = 16'sd5;
        fc1_weights[73][104] = 16'sd-41;
        fc1_weights[73][105] = 16'sd22;
        fc1_weights[73][106] = 16'sd-62;
        fc1_weights[73][107] = 16'sd-42;
        fc1_weights[73][108] = 16'sd-47;
        fc1_weights[73][109] = 16'sd18;
        fc1_weights[73][110] = 16'sd-33;
        fc1_weights[73][111] = 16'sd15;
        fc1_weights[73][112] = 16'sd-3;
        fc1_weights[73][113] = 16'sd3;
        fc1_weights[73][114] = 16'sd45;
        fc1_weights[73][115] = 16'sd63;
        fc1_weights[73][116] = 16'sd-14;
        fc1_weights[73][117] = 16'sd1;
        fc1_weights[73][118] = 16'sd0;
        fc1_weights[73][119] = 16'sd-74;
        fc1_weights[73][120] = 16'sd-31;
        fc1_weights[73][121] = 16'sd-16;
        fc1_weights[73][122] = 16'sd-76;
        fc1_weights[73][123] = 16'sd-69;
        fc1_weights[73][124] = 16'sd-30;
        fc1_weights[73][125] = 16'sd-47;
        fc1_weights[73][126] = 16'sd32;
        fc1_weights[73][127] = 16'sd-10;
        fc1_weights[73][128] = 16'sd-5;
        fc1_weights[73][129] = 16'sd6;
        fc1_weights[73][130] = 16'sd-6;
        fc1_weights[73][131] = 16'sd-41;
        fc1_weights[73][132] = 16'sd-41;
        fc1_weights[73][133] = 16'sd-61;
        fc1_weights[73][134] = 16'sd0;
        fc1_weights[73][135] = 16'sd7;
        fc1_weights[73][136] = 16'sd-4;
        fc1_weights[73][137] = 16'sd-9;
        fc1_weights[73][138] = 16'sd-37;
        fc1_weights[73][139] = 16'sd-32;
        fc1_weights[73][140] = 16'sd-3;
        fc1_weights[73][141] = 16'sd2;
        fc1_weights[73][142] = 16'sd-13;
        fc1_weights[73][143] = 16'sd24;
        fc1_weights[73][144] = 16'sd7;
        fc1_weights[73][145] = 16'sd1;
        fc1_weights[73][146] = 16'sd-27;
        fc1_weights[73][147] = 16'sd-94;
        fc1_weights[73][148] = 16'sd-85;
        fc1_weights[73][149] = 16'sd-3;
        fc1_weights[73][150] = 16'sd-4;
        fc1_weights[73][151] = 16'sd-26;
        fc1_weights[73][152] = 16'sd-16;
        fc1_weights[73][153] = 16'sd-38;
        fc1_weights[73][154] = 16'sd-24;
        fc1_weights[73][155] = 16'sd1;
        fc1_weights[73][156] = 16'sd-58;
        fc1_weights[73][157] = 16'sd-33;
        fc1_weights[73][158] = 16'sd29;
        fc1_weights[73][159] = 16'sd20;
        fc1_weights[73][160] = 16'sd45;
        fc1_weights[73][161] = 16'sd-12;
        fc1_weights[73][162] = 16'sd10;
        fc1_weights[73][163] = 16'sd-73;
        fc1_weights[73][164] = 16'sd-1;
        fc1_weights[73][165] = 16'sd29;
        fc1_weights[73][166] = 16'sd13;
        fc1_weights[73][167] = 16'sd-10;
        fc1_weights[73][168] = 16'sd19;
        fc1_weights[73][169] = 16'sd0;
        fc1_weights[73][170] = 16'sd2;
        fc1_weights[73][171] = 16'sd57;
        fc1_weights[73][172] = 16'sd43;
        fc1_weights[73][173] = 16'sd22;
        fc1_weights[73][174] = 16'sd4;
        fc1_weights[73][175] = 16'sd26;
        fc1_weights[73][176] = 16'sd5;
        fc1_weights[73][177] = 16'sd-45;
        fc1_weights[73][178] = 16'sd-19;
        fc1_weights[73][179] = 16'sd-3;
        fc1_weights[73][180] = 16'sd-30;
        fc1_weights[73][181] = 16'sd1;
        fc1_weights[73][182] = 16'sd0;
        fc1_weights[73][183] = 16'sd25;
        fc1_weights[73][184] = 16'sd53;
        fc1_weights[73][185] = 16'sd19;
        fc1_weights[73][186] = 16'sd41;
        fc1_weights[73][187] = 16'sd52;
        fc1_weights[73][188] = 16'sd57;
        fc1_weights[73][189] = 16'sd59;
        fc1_weights[73][190] = 16'sd21;
        fc1_weights[73][191] = 16'sd20;
        fc1_weights[73][192] = 16'sd25;
        fc1_weights[73][193] = 16'sd44;
        fc1_weights[73][194] = 16'sd25;
        fc1_weights[73][195] = 16'sd1;
        fc1_weights[73][196] = 16'sd-18;
        fc1_weights[73][197] = 16'sd-19;
        fc1_weights[73][198] = 16'sd58;
        fc1_weights[73][199] = 16'sd10;
        fc1_weights[73][200] = 16'sd13;
        fc1_weights[73][201] = 16'sd45;
        fc1_weights[73][202] = 16'sd-28;
        fc1_weights[73][203] = 16'sd-45;
        fc1_weights[73][204] = 16'sd-6;
        fc1_weights[73][205] = 16'sd-25;
        fc1_weights[73][206] = 16'sd-20;
        fc1_weights[73][207] = 16'sd19;
        fc1_weights[74][0] = 16'sd18;
        fc1_weights[74][1] = 16'sd-41;
        fc1_weights[74][2] = 16'sd-6;
        fc1_weights[74][3] = 16'sd-14;
        fc1_weights[74][4] = 16'sd17;
        fc1_weights[74][5] = 16'sd-9;
        fc1_weights[74][6] = 16'sd27;
        fc1_weights[74][7] = 16'sd16;
        fc1_weights[74][8] = 16'sd-36;
        fc1_weights[74][9] = 16'sd18;
        fc1_weights[74][10] = 16'sd-33;
        fc1_weights[74][11] = 16'sd-24;
        fc1_weights[74][12] = 16'sd-70;
        fc1_weights[74][13] = 16'sd-48;
        fc1_weights[74][14] = 16'sd27;
        fc1_weights[74][15] = 16'sd32;
        fc1_weights[74][16] = 16'sd24;
        fc1_weights[74][17] = 16'sd-31;
        fc1_weights[74][18] = 16'sd-29;
        fc1_weights[74][19] = 16'sd-37;
        fc1_weights[74][20] = 16'sd-7;
        fc1_weights[74][21] = 16'sd-8;
        fc1_weights[74][22] = 16'sd-19;
        fc1_weights[74][23] = 16'sd-19;
        fc1_weights[74][24] = 16'sd14;
        fc1_weights[74][25] = 16'sd-6;
        fc1_weights[74][26] = 16'sd11;
        fc1_weights[74][27] = 16'sd12;
        fc1_weights[74][28] = 16'sd4;
        fc1_weights[74][29] = 16'sd-23;
        fc1_weights[74][30] = 16'sd9;
        fc1_weights[74][31] = 16'sd-18;
        fc1_weights[74][32] = 16'sd-20;
        fc1_weights[74][33] = 16'sd1;
        fc1_weights[74][34] = 16'sd-30;
        fc1_weights[74][35] = 16'sd-12;
        fc1_weights[74][36] = 16'sd17;
        fc1_weights[74][37] = 16'sd-71;
        fc1_weights[74][38] = 16'sd-46;
        fc1_weights[74][39] = 16'sd-4;
        fc1_weights[74][40] = 16'sd45;
        fc1_weights[74][41] = 16'sd43;
        fc1_weights[74][42] = 16'sd-35;
        fc1_weights[74][43] = 16'sd-3;
        fc1_weights[74][44] = 16'sd-17;
        fc1_weights[74][45] = 16'sd-50;
        fc1_weights[74][46] = 16'sd7;
        fc1_weights[74][47] = 16'sd2;
        fc1_weights[74][48] = 16'sd3;
        fc1_weights[74][49] = 16'sd-9;
        fc1_weights[74][50] = 16'sd1;
        fc1_weights[74][51] = 16'sd-42;
        fc1_weights[74][52] = 16'sd46;
        fc1_weights[74][53] = 16'sd85;
        fc1_weights[74][54] = 16'sd27;
        fc1_weights[74][55] = 16'sd8;
        fc1_weights[74][56] = 16'sd-20;
        fc1_weights[74][57] = 16'sd6;
        fc1_weights[74][58] = 16'sd35;
        fc1_weights[74][59] = 16'sd-3;
        fc1_weights[74][60] = 16'sd-10;
        fc1_weights[74][61] = 16'sd-7;
        fc1_weights[74][62] = 16'sd10;
        fc1_weights[74][63] = 16'sd-10;
        fc1_weights[74][64] = 16'sd-25;
        fc1_weights[74][65] = 16'sd-29;
        fc1_weights[74][66] = 16'sd3;
        fc1_weights[74][67] = 16'sd-5;
        fc1_weights[74][68] = 16'sd-31;
        fc1_weights[74][69] = 16'sd-34;
        fc1_weights[74][70] = 16'sd-42;
        fc1_weights[74][71] = 16'sd-16;
        fc1_weights[74][72] = 16'sd-1;
        fc1_weights[74][73] = 16'sd-29;
        fc1_weights[74][74] = 16'sd-2;
        fc1_weights[74][75] = 16'sd3;
        fc1_weights[74][76] = 16'sd22;
        fc1_weights[74][77] = 16'sd-39;
        fc1_weights[74][78] = 16'sd40;
        fc1_weights[74][79] = 16'sd69;
        fc1_weights[74][80] = 16'sd-5;
        fc1_weights[74][81] = 16'sd-4;
        fc1_weights[74][82] = 16'sd36;
        fc1_weights[74][83] = 16'sd-17;
        fc1_weights[74][84] = 16'sd-1;
        fc1_weights[74][85] = 16'sd-8;
        fc1_weights[74][86] = 16'sd16;
        fc1_weights[74][87] = 16'sd-22;
        fc1_weights[74][88] = 16'sd-4;
        fc1_weights[74][89] = 16'sd-27;
        fc1_weights[74][90] = 16'sd-1;
        fc1_weights[74][91] = 16'sd6;
        fc1_weights[74][92] = 16'sd4;
        fc1_weights[74][93] = 16'sd-23;
        fc1_weights[74][94] = 16'sd-16;
        fc1_weights[74][95] = 16'sd-17;
        fc1_weights[74][96] = 16'sd-31;
        fc1_weights[74][97] = 16'sd-23;
        fc1_weights[74][98] = 16'sd11;
        fc1_weights[74][99] = 16'sd17;
        fc1_weights[74][100] = 16'sd-9;
        fc1_weights[74][101] = 16'sd-20;
        fc1_weights[74][102] = 16'sd-27;
        fc1_weights[74][103] = 16'sd-46;
        fc1_weights[74][104] = 16'sd63;
        fc1_weights[74][105] = 16'sd22;
        fc1_weights[74][106] = 16'sd26;
        fc1_weights[74][107] = 16'sd13;
        fc1_weights[74][108] = 16'sd22;
        fc1_weights[74][109] = 16'sd-9;
        fc1_weights[74][110] = 16'sd16;
        fc1_weights[74][111] = 16'sd-40;
        fc1_weights[74][112] = 16'sd-2;
        fc1_weights[74][113] = 16'sd11;
        fc1_weights[74][114] = 16'sd-29;
        fc1_weights[74][115] = 16'sd-2;
        fc1_weights[74][116] = 16'sd20;
        fc1_weights[74][117] = 16'sd-11;
        fc1_weights[74][118] = 16'sd-4;
        fc1_weights[74][119] = 16'sd7;
        fc1_weights[74][120] = 16'sd27;
        fc1_weights[74][121] = 16'sd3;
        fc1_weights[74][122] = 16'sd3;
        fc1_weights[74][123] = 16'sd0;
        fc1_weights[74][124] = 16'sd-14;
        fc1_weights[74][125] = 16'sd-19;
        fc1_weights[74][126] = 16'sd-62;
        fc1_weights[74][127] = 16'sd-46;
        fc1_weights[74][128] = 16'sd-1;
        fc1_weights[74][129] = 16'sd-55;
        fc1_weights[74][130] = 16'sd15;
        fc1_weights[74][131] = 16'sd7;
        fc1_weights[74][132] = 16'sd9;
        fc1_weights[74][133] = 16'sd20;
        fc1_weights[74][134] = 16'sd30;
        fc1_weights[74][135] = 16'sd-15;
        fc1_weights[74][136] = 16'sd8;
        fc1_weights[74][137] = 16'sd16;
        fc1_weights[74][138] = 16'sd-18;
        fc1_weights[74][139] = 16'sd54;
        fc1_weights[74][140] = 16'sd49;
        fc1_weights[74][141] = 16'sd0;
        fc1_weights[74][142] = 16'sd32;
        fc1_weights[74][143] = 16'sd-7;
        fc1_weights[74][144] = 16'sd-41;
        fc1_weights[74][145] = 16'sd-37;
        fc1_weights[74][146] = 16'sd-38;
        fc1_weights[74][147] = 16'sd18;
        fc1_weights[74][148] = 16'sd12;
        fc1_weights[74][149] = 16'sd-3;
        fc1_weights[74][150] = 16'sd-22;
        fc1_weights[74][151] = 16'sd6;
        fc1_weights[74][152] = 16'sd19;
        fc1_weights[74][153] = 16'sd3;
        fc1_weights[74][154] = 16'sd5;
        fc1_weights[74][155] = 16'sd-22;
        fc1_weights[74][156] = 16'sd41;
        fc1_weights[74][157] = 16'sd46;
        fc1_weights[74][158] = 16'sd36;
        fc1_weights[74][159] = 16'sd18;
        fc1_weights[74][160] = 16'sd10;
        fc1_weights[74][161] = 16'sd22;
        fc1_weights[74][162] = 16'sd30;
        fc1_weights[74][163] = 16'sd53;
        fc1_weights[74][164] = 16'sd46;
        fc1_weights[74][165] = 16'sd13;
        fc1_weights[74][166] = 16'sd38;
        fc1_weights[74][167] = 16'sd31;
        fc1_weights[74][168] = 16'sd23;
        fc1_weights[74][169] = 16'sd8;
        fc1_weights[74][170] = 16'sd17;
        fc1_weights[74][171] = 16'sd1;
        fc1_weights[74][172] = 16'sd-10;
        fc1_weights[74][173] = 16'sd4;
        fc1_weights[74][174] = 16'sd-16;
        fc1_weights[74][175] = 16'sd-9;
        fc1_weights[74][176] = 16'sd-8;
        fc1_weights[74][177] = 16'sd-1;
        fc1_weights[74][178] = 16'sd-30;
        fc1_weights[74][179] = 16'sd-27;
        fc1_weights[74][180] = 16'sd-17;
        fc1_weights[74][181] = 16'sd-45;
        fc1_weights[74][182] = 16'sd19;
        fc1_weights[74][183] = 16'sd26;
        fc1_weights[74][184] = 16'sd3;
        fc1_weights[74][185] = 16'sd33;
        fc1_weights[74][186] = 16'sd41;
        fc1_weights[74][187] = 16'sd27;
        fc1_weights[74][188] = 16'sd-1;
        fc1_weights[74][189] = 16'sd42;
        fc1_weights[74][190] = 16'sd39;
        fc1_weights[74][191] = 16'sd14;
        fc1_weights[74][192] = 16'sd-21;
        fc1_weights[74][193] = 16'sd-16;
        fc1_weights[74][194] = 16'sd-14;
        fc1_weights[74][195] = 16'sd-8;
        fc1_weights[74][196] = 16'sd-5;
        fc1_weights[74][197] = 16'sd-16;
        fc1_weights[74][198] = 16'sd-45;
        fc1_weights[74][199] = 16'sd13;
        fc1_weights[74][200] = 16'sd-31;
        fc1_weights[74][201] = 16'sd-30;
        fc1_weights[74][202] = 16'sd-21;
        fc1_weights[74][203] = 16'sd17;
        fc1_weights[74][204] = 16'sd-20;
        fc1_weights[74][205] = 16'sd2;
        fc1_weights[74][206] = 16'sd-37;
        fc1_weights[74][207] = 16'sd-34;
        fc1_weights[75][0] = 16'sd-34;
        fc1_weights[75][1] = 16'sd-8;
        fc1_weights[75][2] = 16'sd17;
        fc1_weights[75][3] = 16'sd39;
        fc1_weights[75][4] = 16'sd-10;
        fc1_weights[75][5] = 16'sd34;
        fc1_weights[75][6] = 16'sd-13;
        fc1_weights[75][7] = 16'sd1;
        fc1_weights[75][8] = 16'sd18;
        fc1_weights[75][9] = 16'sd16;
        fc1_weights[75][10] = 16'sd-8;
        fc1_weights[75][11] = 16'sd29;
        fc1_weights[75][12] = 16'sd13;
        fc1_weights[75][13] = 16'sd6;
        fc1_weights[75][14] = 16'sd-8;
        fc1_weights[75][15] = 16'sd19;
        fc1_weights[75][16] = 16'sd5;
        fc1_weights[75][17] = 16'sd-16;
        fc1_weights[75][18] = 16'sd-1;
        fc1_weights[75][19] = 16'sd-10;
        fc1_weights[75][20] = 16'sd-29;
        fc1_weights[75][21] = 16'sd-24;
        fc1_weights[75][22] = 16'sd-1;
        fc1_weights[75][23] = 16'sd53;
        fc1_weights[75][24] = 16'sd-44;
        fc1_weights[75][25] = 16'sd-22;
        fc1_weights[75][26] = 16'sd26;
        fc1_weights[75][27] = 16'sd-2;
        fc1_weights[75][28] = 16'sd45;
        fc1_weights[75][29] = 16'sd68;
        fc1_weights[75][30] = 16'sd57;
        fc1_weights[75][31] = 16'sd70;
        fc1_weights[75][32] = 16'sd14;
        fc1_weights[75][33] = 16'sd-8;
        fc1_weights[75][34] = 16'sd14;
        fc1_weights[75][35] = 16'sd-26;
        fc1_weights[75][36] = 16'sd8;
        fc1_weights[75][37] = 16'sd63;
        fc1_weights[75][38] = 16'sd23;
        fc1_weights[75][39] = 16'sd39;
        fc1_weights[75][40] = 16'sd5;
        fc1_weights[75][41] = 16'sd-23;
        fc1_weights[75][42] = 16'sd10;
        fc1_weights[75][43] = 16'sd-47;
        fc1_weights[75][44] = 16'sd-28;
        fc1_weights[75][45] = 16'sd-52;
        fc1_weights[75][46] = 16'sd-76;
        fc1_weights[75][47] = 16'sd-40;
        fc1_weights[75][48] = 16'sd-33;
        fc1_weights[75][49] = 16'sd-13;
        fc1_weights[75][50] = 16'sd-30;
        fc1_weights[75][51] = 16'sd-14;
        fc1_weights[75][52] = 16'sd85;
        fc1_weights[75][53] = 16'sd-5;
        fc1_weights[75][54] = 16'sd-6;
        fc1_weights[75][55] = 16'sd4;
        fc1_weights[75][56] = 16'sd22;
        fc1_weights[75][57] = 16'sd8;
        fc1_weights[75][58] = 16'sd-5;
        fc1_weights[75][59] = 16'sd18;
        fc1_weights[75][60] = 16'sd11;
        fc1_weights[75][61] = 16'sd17;
        fc1_weights[75][62] = 16'sd-48;
        fc1_weights[75][63] = 16'sd-33;
        fc1_weights[75][64] = 16'sd1;
        fc1_weights[75][65] = 16'sd-12;
        fc1_weights[75][66] = 16'sd32;
        fc1_weights[75][67] = 16'sd-27;
        fc1_weights[75][68] = 16'sd-65;
        fc1_weights[75][69] = 16'sd-14;
        fc1_weights[75][70] = 16'sd-21;
        fc1_weights[75][71] = 16'sd6;
        fc1_weights[75][72] = 16'sd-17;
        fc1_weights[75][73] = 16'sd-3;
        fc1_weights[75][74] = 16'sd2;
        fc1_weights[75][75] = 16'sd-6;
        fc1_weights[75][76] = 16'sd-4;
        fc1_weights[75][77] = 16'sd-10;
        fc1_weights[75][78] = 16'sd41;
        fc1_weights[75][79] = 16'sd42;
        fc1_weights[75][80] = 16'sd13;
        fc1_weights[75][81] = 16'sd3;
        fc1_weights[75][82] = 16'sd8;
        fc1_weights[75][83] = 16'sd57;
        fc1_weights[75][84] = 16'sd-1;
        fc1_weights[75][85] = 16'sd-7;
        fc1_weights[75][86] = 16'sd45;
        fc1_weights[75][87] = 16'sd90;
        fc1_weights[75][88] = 16'sd7;
        fc1_weights[75][89] = 16'sd-11;
        fc1_weights[75][90] = 16'sd20;
        fc1_weights[75][91] = 16'sd7;
        fc1_weights[75][92] = 16'sd26;
        fc1_weights[75][93] = 16'sd-26;
        fc1_weights[75][94] = 16'sd-56;
        fc1_weights[75][95] = 16'sd13;
        fc1_weights[75][96] = 16'sd-14;
        fc1_weights[75][97] = 16'sd31;
        fc1_weights[75][98] = 16'sd6;
        fc1_weights[75][99] = 16'sd-5;
        fc1_weights[75][100] = 16'sd-11;
        fc1_weights[75][101] = 16'sd-14;
        fc1_weights[75][102] = 16'sd-3;
        fc1_weights[75][103] = 16'sd14;
        fc1_weights[75][104] = 16'sd21;
        fc1_weights[75][105] = 16'sd-29;
        fc1_weights[75][106] = 16'sd16;
        fc1_weights[75][107] = 16'sd11;
        fc1_weights[75][108] = 16'sd-9;
        fc1_weights[75][109] = 16'sd18;
        fc1_weights[75][110] = 16'sd-26;
        fc1_weights[75][111] = 16'sd36;
        fc1_weights[75][112] = 16'sd59;
        fc1_weights[75][113] = 16'sd7;
        fc1_weights[75][114] = 16'sd-17;
        fc1_weights[75][115] = 16'sd-2;
        fc1_weights[75][116] = 16'sd6;
        fc1_weights[75][117] = 16'sd3;
        fc1_weights[75][118] = 16'sd16;
        fc1_weights[75][119] = 16'sd21;
        fc1_weights[75][120] = 16'sd1;
        fc1_weights[75][121] = 16'sd30;
        fc1_weights[75][122] = 16'sd38;
        fc1_weights[75][123] = 16'sd79;
        fc1_weights[75][124] = 16'sd40;
        fc1_weights[75][125] = 16'sd-6;
        fc1_weights[75][126] = 16'sd-27;
        fc1_weights[75][127] = 16'sd16;
        fc1_weights[75][128] = 16'sd28;
        fc1_weights[75][129] = 16'sd16;
        fc1_weights[75][130] = 16'sd-25;
        fc1_weights[75][131] = 16'sd-37;
        fc1_weights[75][132] = 16'sd-9;
        fc1_weights[75][133] = 16'sd-11;
        fc1_weights[75][134] = 16'sd-22;
        fc1_weights[75][135] = 16'sd-10;
        fc1_weights[75][136] = 16'sd-42;
        fc1_weights[75][137] = 16'sd-14;
        fc1_weights[75][138] = 16'sd-6;
        fc1_weights[75][139] = 16'sd-4;
        fc1_weights[75][140] = 16'sd-3;
        fc1_weights[75][141] = 16'sd11;
        fc1_weights[75][142] = 16'sd60;
        fc1_weights[75][143] = 16'sd0;
        fc1_weights[75][144] = 16'sd72;
        fc1_weights[75][145] = 16'sd5;
        fc1_weights[75][146] = 16'sd-9;
        fc1_weights[75][147] = 16'sd-4;
        fc1_weights[75][148] = 16'sd51;
        fc1_weights[75][149] = 16'sd-2;
        fc1_weights[75][150] = 16'sd32;
        fc1_weights[75][151] = 16'sd-17;
        fc1_weights[75][152] = 16'sd-21;
        fc1_weights[75][153] = 16'sd-23;
        fc1_weights[75][154] = 16'sd-24;
        fc1_weights[75][155] = 16'sd-2;
        fc1_weights[75][156] = 16'sd-4;
        fc1_weights[75][157] = 16'sd-1;
        fc1_weights[75][158] = 16'sd-42;
        fc1_weights[75][159] = 16'sd-30;
        fc1_weights[75][160] = 16'sd8;
        fc1_weights[75][161] = 16'sd16;
        fc1_weights[75][162] = 16'sd32;
        fc1_weights[75][163] = 16'sd60;
        fc1_weights[75][164] = 16'sd25;
        fc1_weights[75][165] = 16'sd14;
        fc1_weights[75][166] = 16'sd2;
        fc1_weights[75][167] = 16'sd-16;
        fc1_weights[75][168] = 16'sd27;
        fc1_weights[75][169] = 16'sd15;
        fc1_weights[75][170] = 16'sd4;
        fc1_weights[75][171] = 16'sd22;
        fc1_weights[75][172] = 16'sd-19;
        fc1_weights[75][173] = 16'sd-15;
        fc1_weights[75][174] = 16'sd20;
        fc1_weights[75][175] = 16'sd-11;
        fc1_weights[75][176] = 16'sd-16;
        fc1_weights[75][177] = 16'sd29;
        fc1_weights[75][178] = 16'sd-51;
        fc1_weights[75][179] = 16'sd-28;
        fc1_weights[75][180] = 16'sd-4;
        fc1_weights[75][181] = 16'sd-29;
        fc1_weights[75][182] = 16'sd-15;
        fc1_weights[75][183] = 16'sd-21;
        fc1_weights[75][184] = 16'sd-34;
        fc1_weights[75][185] = 16'sd-24;
        fc1_weights[75][186] = 16'sd17;
        fc1_weights[75][187] = 16'sd-3;
        fc1_weights[75][188] = 16'sd2;
        fc1_weights[75][189] = 16'sd28;
        fc1_weights[75][190] = 16'sd-1;
        fc1_weights[75][191] = 16'sd1;
        fc1_weights[75][192] = 16'sd25;
        fc1_weights[75][193] = 16'sd-6;
        fc1_weights[75][194] = 16'sd52;
        fc1_weights[75][195] = 16'sd17;
        fc1_weights[75][196] = 16'sd8;
        fc1_weights[75][197] = 16'sd11;
        fc1_weights[75][198] = 16'sd10;
        fc1_weights[75][199] = 16'sd-7;
        fc1_weights[75][200] = 16'sd-18;
        fc1_weights[75][201] = 16'sd-1;
        fc1_weights[75][202] = 16'sd47;
        fc1_weights[75][203] = 16'sd7;
        fc1_weights[75][204] = 16'sd14;
        fc1_weights[75][205] = 16'sd-39;
        fc1_weights[75][206] = 16'sd15;
        fc1_weights[75][207] = 16'sd-14;
        fc1_weights[76][0] = 16'sd-13;
        fc1_weights[76][1] = 16'sd-27;
        fc1_weights[76][2] = 16'sd-13;
        fc1_weights[76][3] = 16'sd-2;
        fc1_weights[76][4] = 16'sd-18;
        fc1_weights[76][5] = 16'sd-39;
        fc1_weights[76][6] = 16'sd-5;
        fc1_weights[76][7] = 16'sd-48;
        fc1_weights[76][8] = 16'sd-17;
        fc1_weights[76][9] = 16'sd-33;
        fc1_weights[76][10] = 16'sd-7;
        fc1_weights[76][11] = 16'sd1;
        fc1_weights[76][12] = 16'sd-14;
        fc1_weights[76][13] = 16'sd-11;
        fc1_weights[76][14] = 16'sd-21;
        fc1_weights[76][15] = 16'sd37;
        fc1_weights[76][16] = 16'sd20;
        fc1_weights[76][17] = 16'sd29;
        fc1_weights[76][18] = 16'sd12;
        fc1_weights[76][19] = 16'sd8;
        fc1_weights[76][20] = 16'sd-7;
        fc1_weights[76][21] = 16'sd-33;
        fc1_weights[76][22] = 16'sd-74;
        fc1_weights[76][23] = 16'sd-38;
        fc1_weights[76][24] = 16'sd30;
        fc1_weights[76][25] = 16'sd26;
        fc1_weights[76][26] = 16'sd5;
        fc1_weights[76][27] = 16'sd-19;
        fc1_weights[76][28] = 16'sd-39;
        fc1_weights[76][29] = 16'sd4;
        fc1_weights[76][30] = 16'sd13;
        fc1_weights[76][31] = 16'sd5;
        fc1_weights[76][32] = 16'sd11;
        fc1_weights[76][33] = 16'sd-72;
        fc1_weights[76][34] = 16'sd-3;
        fc1_weights[76][35] = 16'sd-8;
        fc1_weights[76][36] = 16'sd33;
        fc1_weights[76][37] = 16'sd27;
        fc1_weights[76][38] = 16'sd3;
        fc1_weights[76][39] = 16'sd-6;
        fc1_weights[76][40] = 16'sd31;
        fc1_weights[76][41] = 16'sd33;
        fc1_weights[76][42] = 16'sd31;
        fc1_weights[76][43] = 16'sd39;
        fc1_weights[76][44] = 16'sd21;
        fc1_weights[76][45] = 16'sd27;
        fc1_weights[76][46] = 16'sd-6;
        fc1_weights[76][47] = 16'sd-25;
        fc1_weights[76][48] = 16'sd-46;
        fc1_weights[76][49] = 16'sd19;
        fc1_weights[76][50] = 16'sd-6;
        fc1_weights[76][51] = 16'sd19;
        fc1_weights[76][52] = 16'sd-36;
        fc1_weights[76][53] = 16'sd21;
        fc1_weights[76][54] = 16'sd21;
        fc1_weights[76][55] = 16'sd-4;
        fc1_weights[76][56] = 16'sd-8;
        fc1_weights[76][57] = 16'sd-13;
        fc1_weights[76][58] = 16'sd-47;
        fc1_weights[76][59] = 16'sd-26;
        fc1_weights[76][60] = 16'sd-4;
        fc1_weights[76][61] = 16'sd-25;
        fc1_weights[76][62] = 16'sd29;
        fc1_weights[76][63] = 16'sd32;
        fc1_weights[76][64] = 16'sd30;
        fc1_weights[76][65] = 16'sd61;
        fc1_weights[76][66] = 16'sd20;
        fc1_weights[76][67] = 16'sd-24;
        fc1_weights[76][68] = 16'sd-6;
        fc1_weights[76][69] = 16'sd3;
        fc1_weights[76][70] = 16'sd-15;
        fc1_weights[76][71] = 16'sd-31;
        fc1_weights[76][72] = 16'sd-1;
        fc1_weights[76][73] = 16'sd-43;
        fc1_weights[76][74] = 16'sd-13;
        fc1_weights[76][75] = 16'sd-19;
        fc1_weights[76][76] = 16'sd-12;
        fc1_weights[76][77] = 16'sd13;
        fc1_weights[76][78] = 16'sd2;
        fc1_weights[76][79] = 16'sd11;
        fc1_weights[76][80] = 16'sd23;
        fc1_weights[76][81] = 16'sd-1;
        fc1_weights[76][82] = 16'sd-41;
        fc1_weights[76][83] = 16'sd-15;
        fc1_weights[76][84] = 16'sd-42;
        fc1_weights[76][85] = 16'sd-44;
        fc1_weights[76][86] = 16'sd-14;
        fc1_weights[76][87] = 16'sd14;
        fc1_weights[76][88] = 16'sd4;
        fc1_weights[76][89] = 16'sd46;
        fc1_weights[76][90] = 16'sd-5;
        fc1_weights[76][91] = 16'sd-5;
        fc1_weights[76][92] = 16'sd53;
        fc1_weights[76][93] = 16'sd19;
        fc1_weights[76][94] = 16'sd10;
        fc1_weights[76][95] = 16'sd6;
        fc1_weights[76][96] = 16'sd2;
        fc1_weights[76][97] = 16'sd17;
        fc1_weights[76][98] = 16'sd-16;
        fc1_weights[76][99] = 16'sd-38;
        fc1_weights[76][100] = 16'sd18;
        fc1_weights[76][101] = 16'sd11;
        fc1_weights[76][102] = 16'sd-11;
        fc1_weights[76][103] = 16'sd-11;
        fc1_weights[76][104] = 16'sd0;
        fc1_weights[76][105] = 16'sd26;
        fc1_weights[76][106] = 16'sd-17;
        fc1_weights[76][107] = 16'sd-4;
        fc1_weights[76][108] = 16'sd18;
        fc1_weights[76][109] = 16'sd16;
        fc1_weights[76][110] = 16'sd-39;
        fc1_weights[76][111] = 16'sd21;
        fc1_weights[76][112] = 16'sd19;
        fc1_weights[76][113] = 16'sd30;
        fc1_weights[76][114] = 16'sd23;
        fc1_weights[76][115] = 16'sd56;
        fc1_weights[76][116] = 16'sd61;
        fc1_weights[76][117] = 16'sd72;
        fc1_weights[76][118] = 16'sd33;
        fc1_weights[76][119] = 16'sd42;
        fc1_weights[76][120] = 16'sd-3;
        fc1_weights[76][121] = 16'sd4;
        fc1_weights[76][122] = 16'sd30;
        fc1_weights[76][123] = 16'sd93;
        fc1_weights[76][124] = 16'sd-9;
        fc1_weights[76][125] = 16'sd5;
        fc1_weights[76][126] = 16'sd12;
        fc1_weights[76][127] = 16'sd28;
        fc1_weights[76][128] = 16'sd11;
        fc1_weights[76][129] = 16'sd-14;
        fc1_weights[76][130] = 16'sd-71;
        fc1_weights[76][131] = 16'sd-55;
        fc1_weights[76][132] = 16'sd-5;
        fc1_weights[76][133] = 16'sd-13;
        fc1_weights[76][134] = 16'sd29;
        fc1_weights[76][135] = 16'sd2;
        fc1_weights[76][136] = 16'sd-48;
        fc1_weights[76][137] = 16'sd-30;
        fc1_weights[76][138] = 16'sd46;
        fc1_weights[76][139] = 16'sd36;
        fc1_weights[76][140] = 16'sd60;
        fc1_weights[76][141] = 16'sd25;
        fc1_weights[76][142] = 16'sd50;
        fc1_weights[76][143] = 16'sd31;
        fc1_weights[76][144] = 16'sd36;
        fc1_weights[76][145] = 16'sd-12;
        fc1_weights[76][146] = 16'sd11;
        fc1_weights[76][147] = 16'sd-16;
        fc1_weights[76][148] = 16'sd35;
        fc1_weights[76][149] = 16'sd55;
        fc1_weights[76][150] = 16'sd-2;
        fc1_weights[76][151] = 16'sd33;
        fc1_weights[76][152] = 16'sd-31;
        fc1_weights[76][153] = 16'sd-12;
        fc1_weights[76][154] = 16'sd-37;
        fc1_weights[76][155] = 16'sd0;
        fc1_weights[76][156] = 16'sd-18;
        fc1_weights[76][157] = 16'sd-9;
        fc1_weights[76][158] = 16'sd1;
        fc1_weights[76][159] = 16'sd15;
        fc1_weights[76][160] = 16'sd-15;
        fc1_weights[76][161] = 16'sd-31;
        fc1_weights[76][162] = 16'sd63;
        fc1_weights[76][163] = 16'sd44;
        fc1_weights[76][164] = 16'sd21;
        fc1_weights[76][165] = 16'sd-21;
        fc1_weights[76][166] = 16'sd4;
        fc1_weights[76][167] = 16'sd19;
        fc1_weights[76][168] = 16'sd50;
        fc1_weights[76][169] = 16'sd-15;
        fc1_weights[76][170] = 16'sd46;
        fc1_weights[76][171] = 16'sd46;
        fc1_weights[76][172] = 16'sd47;
        fc1_weights[76][173] = 16'sd17;
        fc1_weights[76][174] = 16'sd-16;
        fc1_weights[76][175] = 16'sd15;
        fc1_weights[76][176] = 16'sd22;
        fc1_weights[76][177] = 16'sd39;
        fc1_weights[76][178] = 16'sd-31;
        fc1_weights[76][179] = 16'sd-1;
        fc1_weights[76][180] = 16'sd19;
        fc1_weights[76][181] = 16'sd14;
        fc1_weights[76][182] = 16'sd-31;
        fc1_weights[76][183] = 16'sd7;
        fc1_weights[76][184] = 16'sd-18;
        fc1_weights[76][185] = 16'sd25;
        fc1_weights[76][186] = 16'sd41;
        fc1_weights[76][187] = 16'sd39;
        fc1_weights[76][188] = 16'sd61;
        fc1_weights[76][189] = 16'sd32;
        fc1_weights[76][190] = 16'sd0;
        fc1_weights[76][191] = 16'sd13;
        fc1_weights[76][192] = 16'sd-15;
        fc1_weights[76][193] = 16'sd-18;
        fc1_weights[76][194] = 16'sd-13;
        fc1_weights[76][195] = 16'sd2;
        fc1_weights[76][196] = 16'sd14;
        fc1_weights[76][197] = 16'sd78;
        fc1_weights[76][198] = 16'sd3;
        fc1_weights[76][199] = 16'sd10;
        fc1_weights[76][200] = 16'sd15;
        fc1_weights[76][201] = 16'sd-25;
        fc1_weights[76][202] = 16'sd8;
        fc1_weights[76][203] = 16'sd7;
        fc1_weights[76][204] = 16'sd26;
        fc1_weights[76][205] = 16'sd17;
        fc1_weights[76][206] = 16'sd-19;
        fc1_weights[76][207] = 16'sd-10;
        fc1_weights[77][0] = 16'sd-37;
        fc1_weights[77][1] = 16'sd-2;
        fc1_weights[77][2] = 16'sd-50;
        fc1_weights[77][3] = 16'sd-18;
        fc1_weights[77][4] = 16'sd-44;
        fc1_weights[77][5] = 16'sd13;
        fc1_weights[77][6] = 16'sd-71;
        fc1_weights[77][7] = 16'sd-2;
        fc1_weights[77][8] = 16'sd-40;
        fc1_weights[77][9] = 16'sd-20;
        fc1_weights[77][10] = 16'sd-5;
        fc1_weights[77][11] = 16'sd59;
        fc1_weights[77][12] = 16'sd92;
        fc1_weights[77][13] = 16'sd27;
        fc1_weights[77][14] = 16'sd11;
        fc1_weights[77][15] = 16'sd16;
        fc1_weights[77][16] = 16'sd-28;
        fc1_weights[77][17] = 16'sd-70;
        fc1_weights[77][18] = 16'sd-31;
        fc1_weights[77][19] = 16'sd-5;
        fc1_weights[77][20] = 16'sd-5;
        fc1_weights[77][21] = 16'sd-18;
        fc1_weights[77][22] = 16'sd-54;
        fc1_weights[77][23] = 16'sd-27;
        fc1_weights[77][24] = 16'sd38;
        fc1_weights[77][25] = 16'sd-32;
        fc1_weights[77][26] = 16'sd-66;
        fc1_weights[77][27] = 16'sd-82;
        fc1_weights[77][28] = 16'sd-3;
        fc1_weights[77][29] = 16'sd71;
        fc1_weights[77][30] = 16'sd-35;
        fc1_weights[77][31] = 16'sd-19;
        fc1_weights[77][32] = 16'sd-7;
        fc1_weights[77][33] = 16'sd-107;
        fc1_weights[77][34] = 16'sd-36;
        fc1_weights[77][35] = 16'sd-63;
        fc1_weights[77][36] = 16'sd61;
        fc1_weights[77][37] = 16'sd-15;
        fc1_weights[77][38] = 16'sd28;
        fc1_weights[77][39] = 16'sd1;
        fc1_weights[77][40] = 16'sd57;
        fc1_weights[77][41] = 16'sd-21;
        fc1_weights[77][42] = 16'sd47;
        fc1_weights[77][43] = 16'sd-65;
        fc1_weights[77][44] = 16'sd-22;
        fc1_weights[77][45] = 16'sd89;
        fc1_weights[77][46] = 16'sd27;
        fc1_weights[77][47] = 16'sd-6;
        fc1_weights[77][48] = 16'sd-69;
        fc1_weights[77][49] = 16'sd-48;
        fc1_weights[77][50] = 16'sd6;
        fc1_weights[77][51] = 16'sd31;
        fc1_weights[77][52] = 16'sd33;
        fc1_weights[77][53] = 16'sd24;
        fc1_weights[77][54] = 16'sd-9;
        fc1_weights[77][55] = 16'sd32;
        fc1_weights[77][56] = 16'sd71;
        fc1_weights[77][57] = 16'sd24;
        fc1_weights[77][58] = 16'sd-31;
        fc1_weights[77][59] = 16'sd-45;
        fc1_weights[77][60] = 16'sd77;
        fc1_weights[77][61] = 16'sd21;
        fc1_weights[77][62] = 16'sd-34;
        fc1_weights[77][63] = 16'sd-16;
        fc1_weights[77][64] = 16'sd151;
        fc1_weights[77][65] = 16'sd-2;
        fc1_weights[77][66] = 16'sd40;
        fc1_weights[77][67] = 16'sd-5;
        fc1_weights[77][68] = 16'sd-83;
        fc1_weights[77][69] = 16'sd10;
        fc1_weights[77][70] = 16'sd20;
        fc1_weights[77][71] = 16'sd122;
        fc1_weights[77][72] = 16'sd105;
        fc1_weights[77][73] = 16'sd67;
        fc1_weights[77][74] = 16'sd40;
        fc1_weights[77][75] = 16'sd-38;
        fc1_weights[77][76] = 16'sd-18;
        fc1_weights[77][77] = 16'sd46;
        fc1_weights[77][78] = 16'sd-26;
        fc1_weights[77][79] = 16'sd52;
        fc1_weights[77][80] = 16'sd-31;
        fc1_weights[77][81] = 16'sd59;
        fc1_weights[77][82] = 16'sd48;
        fc1_weights[77][83] = 16'sd70;
        fc1_weights[77][84] = 16'sd51;
        fc1_weights[77][85] = 16'sd2;
        fc1_weights[77][86] = 16'sd28;
        fc1_weights[77][87] = 16'sd99;
        fc1_weights[77][88] = 16'sd48;
        fc1_weights[77][89] = 16'sd-43;
        fc1_weights[77][90] = 16'sd103;
        fc1_weights[77][91] = 16'sd117;
        fc1_weights[77][92] = 16'sd62;
        fc1_weights[77][93] = 16'sd-44;
        fc1_weights[77][94] = 16'sd-113;
        fc1_weights[77][95] = 16'sd39;
        fc1_weights[77][96] = 16'sd-37;
        fc1_weights[77][97] = 16'sd-12;
        fc1_weights[77][98] = 16'sd35;
        fc1_weights[77][99] = 16'sd-64;
        fc1_weights[77][100] = 16'sd32;
        fc1_weights[77][101] = 16'sd3;
        fc1_weights[77][102] = 16'sd-57;
        fc1_weights[77][103] = 16'sd-19;
        fc1_weights[77][104] = 16'sd80;
        fc1_weights[77][105] = 16'sd-32;
        fc1_weights[77][106] = 16'sd63;
        fc1_weights[77][107] = 16'sd17;
        fc1_weights[77][108] = 16'sd-10;
        fc1_weights[77][109] = 16'sd52;
        fc1_weights[77][110] = 16'sd-33;
        fc1_weights[77][111] = 16'sd-8;
        fc1_weights[77][112] = 16'sd70;
        fc1_weights[77][113] = 16'sd-15;
        fc1_weights[77][114] = 16'sd75;
        fc1_weights[77][115] = 16'sd82;
        fc1_weights[77][116] = 16'sd108;
        fc1_weights[77][117] = 16'sd70;
        fc1_weights[77][118] = 16'sd25;
        fc1_weights[77][119] = 16'sd-49;
        fc1_weights[77][120] = 16'sd-12;
        fc1_weights[77][121] = 16'sd42;
        fc1_weights[77][122] = 16'sd36;
        fc1_weights[77][123] = 16'sd-32;
        fc1_weights[77][124] = 16'sd-19;
        fc1_weights[77][125] = 16'sd25;
        fc1_weights[77][126] = 16'sd26;
        fc1_weights[77][127] = 16'sd67;
        fc1_weights[77][128] = 16'sd18;
        fc1_weights[77][129] = 16'sd49;
        fc1_weights[77][130] = 16'sd-60;
        fc1_weights[77][131] = 16'sd-23;
        fc1_weights[77][132] = 16'sd6;
        fc1_weights[77][133] = 16'sd-25;
        fc1_weights[77][134] = 16'sd-5;
        fc1_weights[77][135] = 16'sd28;
        fc1_weights[77][136] = 16'sd44;
        fc1_weights[77][137] = 16'sd25;
        fc1_weights[77][138] = 16'sd74;
        fc1_weights[77][139] = 16'sd-97;
        fc1_weights[77][140] = 16'sd-80;
        fc1_weights[77][141] = 16'sd76;
        fc1_weights[77][142] = 16'sd15;
        fc1_weights[77][143] = 16'sd17;
        fc1_weights[77][144] = 16'sd36;
        fc1_weights[77][145] = 16'sd38;
        fc1_weights[77][146] = 16'sd-4;
        fc1_weights[77][147] = 16'sd-46;
        fc1_weights[77][148] = 16'sd-27;
        fc1_weights[77][149] = 16'sd10;
        fc1_weights[77][150] = 16'sd41;
        fc1_weights[77][151] = 16'sd82;
        fc1_weights[77][152] = 16'sd8;
        fc1_weights[77][153] = 16'sd-13;
        fc1_weights[77][154] = 16'sd19;
        fc1_weights[77][155] = 16'sd54;
        fc1_weights[77][156] = 16'sd-75;
        fc1_weights[77][157] = 16'sd-109;
        fc1_weights[77][158] = 16'sd-56;
        fc1_weights[77][159] = 16'sd11;
        fc1_weights[77][160] = 16'sd-40;
        fc1_weights[77][161] = 16'sd28;
        fc1_weights[77][162] = 16'sd39;
        fc1_weights[77][163] = 16'sd-35;
        fc1_weights[77][164] = 16'sd-59;
        fc1_weights[77][165] = 16'sd-93;
        fc1_weights[77][166] = 16'sd-58;
        fc1_weights[77][167] = 16'sd-63;
        fc1_weights[77][168] = 16'sd-14;
        fc1_weights[77][169] = 16'sd23;
        fc1_weights[77][170] = 16'sd69;
        fc1_weights[77][171] = 16'sd-70;
        fc1_weights[77][172] = 16'sd9;
        fc1_weights[77][173] = 16'sd-49;
        fc1_weights[77][174] = 16'sd-23;
        fc1_weights[77][175] = 16'sd-25;
        fc1_weights[77][176] = 16'sd-27;
        fc1_weights[77][177] = 16'sd28;
        fc1_weights[77][178] = 16'sd49;
        fc1_weights[77][179] = 16'sd0;
        fc1_weights[77][180] = 16'sd3;
        fc1_weights[77][181] = 16'sd12;
        fc1_weights[77][182] = 16'sd46;
        fc1_weights[77][183] = 16'sd-10;
        fc1_weights[77][184] = 16'sd5;
        fc1_weights[77][185] = 16'sd7;
        fc1_weights[77][186] = 16'sd-32;
        fc1_weights[77][187] = 16'sd-50;
        fc1_weights[77][188] = 16'sd-23;
        fc1_weights[77][189] = 16'sd-13;
        fc1_weights[77][190] = 16'sd-1;
        fc1_weights[77][191] = 16'sd-21;
        fc1_weights[77][192] = 16'sd52;
        fc1_weights[77][193] = 16'sd15;
        fc1_weights[77][194] = 16'sd-40;
        fc1_weights[77][195] = 16'sd13;
        fc1_weights[77][196] = 16'sd-1;
        fc1_weights[77][197] = 16'sd45;
        fc1_weights[77][198] = 16'sd-85;
        fc1_weights[77][199] = 16'sd-9;
        fc1_weights[77][200] = 16'sd51;
        fc1_weights[77][201] = 16'sd-11;
        fc1_weights[77][202] = 16'sd-98;
        fc1_weights[77][203] = 16'sd-3;
        fc1_weights[77][204] = 16'sd17;
        fc1_weights[77][205] = 16'sd-41;
        fc1_weights[77][206] = 16'sd49;
        fc1_weights[77][207] = 16'sd32;
        fc1_weights[78][0] = 16'sd-11;
        fc1_weights[78][1] = 16'sd36;
        fc1_weights[78][2] = 16'sd14;
        fc1_weights[78][3] = 16'sd-6;
        fc1_weights[78][4] = 16'sd-13;
        fc1_weights[78][5] = 16'sd4;
        fc1_weights[78][6] = 16'sd-2;
        fc1_weights[78][7] = 16'sd-14;
        fc1_weights[78][8] = 16'sd-17;
        fc1_weights[78][9] = 16'sd-6;
        fc1_weights[78][10] = 16'sd-1;
        fc1_weights[78][11] = 16'sd6;
        fc1_weights[78][12] = 16'sd-31;
        fc1_weights[78][13] = 16'sd-39;
        fc1_weights[78][14] = 16'sd-63;
        fc1_weights[78][15] = 16'sd-48;
        fc1_weights[78][16] = 16'sd-12;
        fc1_weights[78][17] = 16'sd-32;
        fc1_weights[78][18] = 16'sd-24;
        fc1_weights[78][19] = 16'sd0;
        fc1_weights[78][20] = 16'sd-1;
        fc1_weights[78][21] = 16'sd-19;
        fc1_weights[78][22] = 16'sd0;
        fc1_weights[78][23] = 16'sd32;
        fc1_weights[78][24] = 16'sd11;
        fc1_weights[78][25] = 16'sd-5;
        fc1_weights[78][26] = 16'sd-37;
        fc1_weights[78][27] = 16'sd-4;
        fc1_weights[78][28] = 16'sd12;
        fc1_weights[78][29] = 16'sd-16;
        fc1_weights[78][30] = 16'sd-11;
        fc1_weights[78][31] = 16'sd19;
        fc1_weights[78][32] = 16'sd29;
        fc1_weights[78][33] = 16'sd49;
        fc1_weights[78][34] = 16'sd17;
        fc1_weights[78][35] = 16'sd16;
        fc1_weights[78][36] = 16'sd10;
        fc1_weights[78][37] = 16'sd-11;
        fc1_weights[78][38] = 16'sd-9;
        fc1_weights[78][39] = 16'sd-32;
        fc1_weights[78][40] = 16'sd-6;
        fc1_weights[78][41] = 16'sd-32;
        fc1_weights[78][42] = 16'sd-40;
        fc1_weights[78][43] = 16'sd5;
        fc1_weights[78][44] = 16'sd-7;
        fc1_weights[78][45] = 16'sd-22;
        fc1_weights[78][46] = 16'sd-4;
        fc1_weights[78][47] = 16'sd4;
        fc1_weights[78][48] = 16'sd-35;
        fc1_weights[78][49] = 16'sd-19;
        fc1_weights[78][50] = 16'sd-3;
        fc1_weights[78][51] = 16'sd-36;
        fc1_weights[78][52] = 16'sd-30;
        fc1_weights[78][53] = 16'sd-2;
        fc1_weights[78][54] = 16'sd32;
        fc1_weights[78][55] = 16'sd33;
        fc1_weights[78][56] = 16'sd3;
        fc1_weights[78][57] = 16'sd13;
        fc1_weights[78][58] = 16'sd19;
        fc1_weights[78][59] = 16'sd14;
        fc1_weights[78][60] = 16'sd-19;
        fc1_weights[78][61] = 16'sd-24;
        fc1_weights[78][62] = 16'sd20;
        fc1_weights[78][63] = 16'sd3;
        fc1_weights[78][64] = 16'sd24;
        fc1_weights[78][65] = 16'sd-22;
        fc1_weights[78][66] = 16'sd-32;
        fc1_weights[78][67] = 16'sd-18;
        fc1_weights[78][68] = 16'sd-10;
        fc1_weights[78][69] = 16'sd20;
        fc1_weights[78][70] = 16'sd-5;
        fc1_weights[78][71] = 16'sd7;
        fc1_weights[78][72] = 16'sd52;
        fc1_weights[78][73] = 16'sd-22;
        fc1_weights[78][74] = 16'sd-51;
        fc1_weights[78][75] = 16'sd40;
        fc1_weights[78][76] = 16'sd11;
        fc1_weights[78][77] = 16'sd6;
        fc1_weights[78][78] = 16'sd-11;
        fc1_weights[78][79] = 16'sd-7;
        fc1_weights[78][80] = 16'sd34;
        fc1_weights[78][81] = 16'sd3;
        fc1_weights[78][82] = 16'sd-2;
        fc1_weights[78][83] = 16'sd-12;
        fc1_weights[78][84] = 16'sd17;
        fc1_weights[78][85] = 16'sd35;
        fc1_weights[78][86] = 16'sd33;
        fc1_weights[78][87] = 16'sd18;
        fc1_weights[78][88] = 16'sd-22;
        fc1_weights[78][89] = 16'sd35;
        fc1_weights[78][90] = 16'sd36;
        fc1_weights[78][91] = 16'sd-8;
        fc1_weights[78][92] = 16'sd-3;
        fc1_weights[78][93] = 16'sd8;
        fc1_weights[78][94] = 16'sd35;
        fc1_weights[78][95] = 16'sd2;
        fc1_weights[78][96] = 16'sd-8;
        fc1_weights[78][97] = 16'sd-52;
        fc1_weights[78][98] = 16'sd10;
        fc1_weights[78][99] = 16'sd9;
        fc1_weights[78][100] = 16'sd-21;
        fc1_weights[78][101] = 16'sd19;
        fc1_weights[78][102] = 16'sd63;
        fc1_weights[78][103] = 16'sd17;
        fc1_weights[78][104] = 16'sd-46;
        fc1_weights[78][105] = 16'sd-24;
        fc1_weights[78][106] = 16'sd-3;
        fc1_weights[78][107] = 16'sd-16;
        fc1_weights[78][108] = 16'sd-3;
        fc1_weights[78][109] = 16'sd-16;
        fc1_weights[78][110] = 16'sd34;
        fc1_weights[78][111] = 16'sd46;
        fc1_weights[78][112] = 16'sd-2;
        fc1_weights[78][113] = 16'sd27;
        fc1_weights[78][114] = 16'sd-4;
        fc1_weights[78][115] = 16'sd-31;
        fc1_weights[78][116] = 16'sd-11;
        fc1_weights[78][117] = 16'sd10;
        fc1_weights[78][118] = 16'sd18;
        fc1_weights[78][119] = 16'sd11;
        fc1_weights[78][120] = 16'sd-1;
        fc1_weights[78][121] = 16'sd1;
        fc1_weights[78][122] = 16'sd5;
        fc1_weights[78][123] = 16'sd-16;
        fc1_weights[78][124] = 16'sd28;
        fc1_weights[78][125] = 16'sd41;
        fc1_weights[78][126] = 16'sd-21;
        fc1_weights[78][127] = 16'sd37;
        fc1_weights[78][128] = 16'sd25;
        fc1_weights[78][129] = 16'sd14;
        fc1_weights[78][130] = 16'sd6;
        fc1_weights[78][131] = 16'sd-28;
        fc1_weights[78][132] = 16'sd7;
        fc1_weights[78][133] = 16'sd-44;
        fc1_weights[78][134] = 16'sd-21;
        fc1_weights[78][135] = 16'sd-2;
        fc1_weights[78][136] = 16'sd-5;
        fc1_weights[78][137] = 16'sd-6;
        fc1_weights[78][138] = 16'sd-45;
        fc1_weights[78][139] = 16'sd27;
        fc1_weights[78][140] = 16'sd-20;
        fc1_weights[78][141] = 16'sd-45;
        fc1_weights[78][142] = 16'sd-14;
        fc1_weights[78][143] = 16'sd-2;
        fc1_weights[78][144] = 16'sd-24;
        fc1_weights[78][145] = 16'sd-38;
        fc1_weights[78][146] = 16'sd-12;
        fc1_weights[78][147] = 16'sd1;
        fc1_weights[78][148] = 16'sd-9;
        fc1_weights[78][149] = 16'sd3;
        fc1_weights[78][150] = 16'sd3;
        fc1_weights[78][151] = 16'sd-2;
        fc1_weights[78][152] = 16'sd30;
        fc1_weights[78][153] = 16'sd39;
        fc1_weights[78][154] = 16'sd48;
        fc1_weights[78][155] = 16'sd32;
        fc1_weights[78][156] = 16'sd8;
        fc1_weights[78][157] = 16'sd0;
        fc1_weights[78][158] = 16'sd16;
        fc1_weights[78][159] = 16'sd-10;
        fc1_weights[78][160] = 16'sd-25;
        fc1_weights[78][161] = 16'sd8;
        fc1_weights[78][162] = 16'sd-5;
        fc1_weights[78][163] = 16'sd20;
        fc1_weights[78][164] = 16'sd25;
        fc1_weights[78][165] = 16'sd7;
        fc1_weights[78][166] = 16'sd-5;
        fc1_weights[78][167] = 16'sd-4;
        fc1_weights[78][168] = 16'sd-12;
        fc1_weights[78][169] = 16'sd-16;
        fc1_weights[78][170] = 16'sd-9;
        fc1_weights[78][171] = 16'sd19;
        fc1_weights[78][172] = 16'sd14;
        fc1_weights[78][173] = 16'sd4;
        fc1_weights[78][174] = 16'sd14;
        fc1_weights[78][175] = 16'sd10;
        fc1_weights[78][176] = 16'sd50;
        fc1_weights[78][177] = 16'sd-3;
        fc1_weights[78][178] = 16'sd-8;
        fc1_weights[78][179] = 16'sd12;
        fc1_weights[78][180] = 16'sd6;
        fc1_weights[78][181] = 16'sd7;
        fc1_weights[78][182] = 16'sd-3;
        fc1_weights[78][183] = 16'sd-7;
        fc1_weights[78][184] = 16'sd-6;
        fc1_weights[78][185] = 16'sd-21;
        fc1_weights[78][186] = 16'sd-23;
        fc1_weights[78][187] = 16'sd2;
        fc1_weights[78][188] = 16'sd-10;
        fc1_weights[78][189] = 16'sd-10;
        fc1_weights[78][190] = 16'sd-9;
        fc1_weights[78][191] = 16'sd-11;
        fc1_weights[78][192] = 16'sd-14;
        fc1_weights[78][193] = 16'sd-14;
        fc1_weights[78][194] = 16'sd-1;
        fc1_weights[78][195] = 16'sd-27;
        fc1_weights[78][196] = 16'sd3;
        fc1_weights[78][197] = 16'sd7;
        fc1_weights[78][198] = 16'sd51;
        fc1_weights[78][199] = 16'sd21;
        fc1_weights[78][200] = 16'sd15;
        fc1_weights[78][201] = 16'sd8;
        fc1_weights[78][202] = 16'sd12;
        fc1_weights[78][203] = 16'sd7;
        fc1_weights[78][204] = 16'sd19;
        fc1_weights[78][205] = 16'sd-16;
        fc1_weights[78][206] = 16'sd-5;
        fc1_weights[78][207] = 16'sd1;
        fc1_weights[79][0] = 16'sd-31;
        fc1_weights[79][1] = 16'sd-2;
        fc1_weights[79][2] = 16'sd-22;
        fc1_weights[79][3] = 16'sd42;
        fc1_weights[79][4] = 16'sd-21;
        fc1_weights[79][5] = 16'sd-18;
        fc1_weights[79][6] = 16'sd-61;
        fc1_weights[79][7] = 16'sd1;
        fc1_weights[79][8] = 16'sd40;
        fc1_weights[79][9] = 16'sd21;
        fc1_weights[79][10] = 16'sd1;
        fc1_weights[79][11] = 16'sd70;
        fc1_weights[79][12] = 16'sd91;
        fc1_weights[79][13] = 16'sd104;
        fc1_weights[79][14] = 16'sd61;
        fc1_weights[79][15] = 16'sd44;
        fc1_weights[79][16] = 16'sd9;
        fc1_weights[79][17] = 16'sd-13;
        fc1_weights[79][18] = 16'sd17;
        fc1_weights[79][19] = 16'sd-5;
        fc1_weights[79][20] = 16'sd9;
        fc1_weights[79][21] = 16'sd40;
        fc1_weights[79][22] = 16'sd-1;
        fc1_weights[79][23] = 16'sd-45;
        fc1_weights[79][24] = 16'sd-19;
        fc1_weights[79][25] = 16'sd-16;
        fc1_weights[79][26] = 16'sd14;
        fc1_weights[79][27] = 16'sd-33;
        fc1_weights[79][28] = 16'sd42;
        fc1_weights[79][29] = 16'sd2;
        fc1_weights[79][30] = 16'sd-39;
        fc1_weights[79][31] = 16'sd-82;
        fc1_weights[79][32] = 16'sd-11;
        fc1_weights[79][33] = 16'sd50;
        fc1_weights[79][34] = 16'sd-3;
        fc1_weights[79][35] = 16'sd-5;
        fc1_weights[79][36] = 16'sd0;
        fc1_weights[79][37] = 16'sd-29;
        fc1_weights[79][38] = 16'sd4;
        fc1_weights[79][39] = 16'sd37;
        fc1_weights[79][40] = 16'sd-7;
        fc1_weights[79][41] = 16'sd32;
        fc1_weights[79][42] = 16'sd44;
        fc1_weights[79][43] = 16'sd43;
        fc1_weights[79][44] = 16'sd32;
        fc1_weights[79][45] = 16'sd69;
        fc1_weights[79][46] = 16'sd35;
        fc1_weights[79][47] = 16'sd79;
        fc1_weights[79][48] = 16'sd13;
        fc1_weights[79][49] = 16'sd-23;
        fc1_weights[79][50] = 16'sd42;
        fc1_weights[79][51] = 16'sd35;
        fc1_weights[79][52] = 16'sd-10;
        fc1_weights[79][53] = 16'sd17;
        fc1_weights[79][54] = 16'sd6;
        fc1_weights[79][55] = 16'sd-6;
        fc1_weights[79][56] = 16'sd-56;
        fc1_weights[79][57] = 16'sd-89;
        fc1_weights[79][58] = 16'sd-21;
        fc1_weights[79][59] = 16'sd-45;
        fc1_weights[79][60] = 16'sd-42;
        fc1_weights[79][61] = 16'sd-29;
        fc1_weights[79][62] = 16'sd52;
        fc1_weights[79][63] = 16'sd33;
        fc1_weights[79][64] = 16'sd-4;
        fc1_weights[79][65] = 16'sd60;
        fc1_weights[79][66] = 16'sd-23;
        fc1_weights[79][67] = 16'sd50;
        fc1_weights[79][68] = 16'sd20;
        fc1_weights[79][69] = 16'sd39;
        fc1_weights[79][70] = 16'sd38;
        fc1_weights[79][71] = 16'sd-1;
        fc1_weights[79][72] = 16'sd-10;
        fc1_weights[79][73] = 16'sd8;
        fc1_weights[79][74] = 16'sd-36;
        fc1_weights[79][75] = 16'sd23;
        fc1_weights[79][76] = 16'sd5;
        fc1_weights[79][77] = 16'sd51;
        fc1_weights[79][78] = 16'sd-32;
        fc1_weights[79][79] = 16'sd-25;
        fc1_weights[79][80] = 16'sd-31;
        fc1_weights[79][81] = 16'sd-32;
        fc1_weights[79][82] = 16'sd-15;
        fc1_weights[79][83] = 16'sd13;
        fc1_weights[79][84] = 16'sd3;
        fc1_weights[79][85] = 16'sd-6;
        fc1_weights[79][86] = 16'sd-20;
        fc1_weights[79][87] = 16'sd-54;
        fc1_weights[79][88] = 16'sd-11;
        fc1_weights[79][89] = 16'sd-4;
        fc1_weights[79][90] = 16'sd-22;
        fc1_weights[79][91] = 16'sd11;
        fc1_weights[79][92] = 16'sd42;
        fc1_weights[79][93] = 16'sd52;
        fc1_weights[79][94] = 16'sd38;
        fc1_weights[79][95] = 16'sd5;
        fc1_weights[79][96] = 16'sd47;
        fc1_weights[79][97] = 16'sd4;
        fc1_weights[79][98] = 16'sd-3;
        fc1_weights[79][99] = 16'sd5;
        fc1_weights[79][100] = 16'sd-20;
        fc1_weights[79][101] = 16'sd33;
        fc1_weights[79][102] = 16'sd55;
        fc1_weights[79][103] = 16'sd37;
        fc1_weights[79][104] = 16'sd-19;
        fc1_weights[79][105] = 16'sd-2;
        fc1_weights[79][106] = 16'sd33;
        fc1_weights[79][107] = 16'sd-8;
        fc1_weights[79][108] = 16'sd-5;
        fc1_weights[79][109] = 16'sd-27;
        fc1_weights[79][110] = 16'sd-13;
        fc1_weights[79][111] = 16'sd19;
        fc1_weights[79][112] = 16'sd-53;
        fc1_weights[79][113] = 16'sd-34;
        fc1_weights[79][114] = 16'sd7;
        fc1_weights[79][115] = 16'sd1;
        fc1_weights[79][116] = 16'sd-18;
        fc1_weights[79][117] = 16'sd-25;
        fc1_weights[79][118] = 16'sd-24;
        fc1_weights[79][119] = 16'sd5;
        fc1_weights[79][120] = 16'sd0;
        fc1_weights[79][121] = 16'sd-27;
        fc1_weights[79][122] = 16'sd-6;
        fc1_weights[79][123] = 16'sd-27;
        fc1_weights[79][124] = 16'sd12;
        fc1_weights[79][125] = 16'sd-12;
        fc1_weights[79][126] = 16'sd15;
        fc1_weights[79][127] = 16'sd-2;
        fc1_weights[79][128] = 16'sd6;
        fc1_weights[79][129] = 16'sd24;
        fc1_weights[79][130] = 16'sd2;
        fc1_weights[79][131] = 16'sd-34;
        fc1_weights[79][132] = 16'sd-29;
        fc1_weights[79][133] = 16'sd10;
        fc1_weights[79][134] = 16'sd2;
        fc1_weights[79][135] = 16'sd15;
        fc1_weights[79][136] = 16'sd-18;
        fc1_weights[79][137] = 16'sd8;
        fc1_weights[79][138] = 16'sd-37;
        fc1_weights[79][139] = 16'sd-49;
        fc1_weights[79][140] = 16'sd-25;
        fc1_weights[79][141] = 16'sd27;
        fc1_weights[79][142] = 16'sd-50;
        fc1_weights[79][143] = 16'sd-29;
        fc1_weights[79][144] = 16'sd-42;
        fc1_weights[79][145] = 16'sd16;
        fc1_weights[79][146] = 16'sd-34;
        fc1_weights[79][147] = 16'sd-42;
        fc1_weights[79][148] = 16'sd-22;
        fc1_weights[79][149] = 16'sd24;
        fc1_weights[79][150] = 16'sd12;
        fc1_weights[79][151] = 16'sd10;
        fc1_weights[79][152] = 16'sd21;
        fc1_weights[79][153] = 16'sd6;
        fc1_weights[79][154] = 16'sd19;
        fc1_weights[79][155] = 16'sd-57;
        fc1_weights[79][156] = 16'sd10;
        fc1_weights[79][157] = 16'sd20;
        fc1_weights[79][158] = 16'sd7;
        fc1_weights[79][159] = 16'sd30;
        fc1_weights[79][160] = 16'sd25;
        fc1_weights[79][161] = 16'sd38;
        fc1_weights[79][162] = 16'sd-4;
        fc1_weights[79][163] = 16'sd24;
        fc1_weights[79][164] = 16'sd-16;
        fc1_weights[79][165] = 16'sd-39;
        fc1_weights[79][166] = 16'sd-31;
        fc1_weights[79][167] = 16'sd-5;
        fc1_weights[79][168] = 16'sd-1;
        fc1_weights[79][169] = 16'sd-10;
        fc1_weights[79][170] = 16'sd-16;
        fc1_weights[79][171] = 16'sd22;
        fc1_weights[79][172] = 16'sd-2;
        fc1_weights[79][173] = 16'sd-10;
        fc1_weights[79][174] = 16'sd-14;
        fc1_weights[79][175] = 16'sd4;
        fc1_weights[79][176] = 16'sd-15;
        fc1_weights[79][177] = 16'sd-16;
        fc1_weights[79][178] = 16'sd4;
        fc1_weights[79][179] = 16'sd-42;
        fc1_weights[79][180] = 16'sd0;
        fc1_weights[79][181] = 16'sd-15;
        fc1_weights[79][182] = 16'sd29;
        fc1_weights[79][183] = 16'sd16;
        fc1_weights[79][184] = 16'sd27;
        fc1_weights[79][185] = 16'sd7;
        fc1_weights[79][186] = 16'sd53;
        fc1_weights[79][187] = 16'sd2;
        fc1_weights[79][188] = 16'sd33;
        fc1_weights[79][189] = 16'sd16;
        fc1_weights[79][190] = 16'sd-59;
        fc1_weights[79][191] = 16'sd-62;
        fc1_weights[79][192] = 16'sd-38;
        fc1_weights[79][193] = 16'sd-20;
        fc1_weights[79][194] = 16'sd-13;
        fc1_weights[79][195] = 16'sd15;
        fc1_weights[79][196] = 16'sd0;
        fc1_weights[79][197] = 16'sd-52;
        fc1_weights[79][198] = 16'sd-17;
        fc1_weights[79][199] = 16'sd-23;
        fc1_weights[79][200] = 16'sd-31;
        fc1_weights[79][201] = 16'sd0;
        fc1_weights[79][202] = 16'sd1;
        fc1_weights[79][203] = 16'sd-61;
        fc1_weights[79][204] = 16'sd-35;
        fc1_weights[79][205] = 16'sd19;
        fc1_weights[79][206] = 16'sd17;
        fc1_weights[79][207] = 16'sd27;
        fc1_weights[80][0] = 16'sd13;
        fc1_weights[80][1] = 16'sd-44;
        fc1_weights[80][2] = 16'sd-14;
        fc1_weights[80][3] = 16'sd-25;
        fc1_weights[80][4] = 16'sd-2;
        fc1_weights[80][5] = 16'sd-39;
        fc1_weights[80][6] = 16'sd-21;
        fc1_weights[80][7] = 16'sd-46;
        fc1_weights[80][8] = 16'sd1;
        fc1_weights[80][9] = 16'sd-1;
        fc1_weights[80][10] = 16'sd-63;
        fc1_weights[80][11] = 16'sd-18;
        fc1_weights[80][12] = 16'sd-17;
        fc1_weights[80][13] = 16'sd-2;
        fc1_weights[80][14] = 16'sd-47;
        fc1_weights[80][15] = 16'sd-49;
        fc1_weights[80][16] = 16'sd-21;
        fc1_weights[80][17] = 16'sd27;
        fc1_weights[80][18] = 16'sd42;
        fc1_weights[80][19] = 16'sd96;
        fc1_weights[80][20] = 16'sd57;
        fc1_weights[80][21] = 16'sd12;
        fc1_weights[80][22] = 16'sd-36;
        fc1_weights[80][23] = 16'sd-2;
        fc1_weights[80][24] = 16'sd-24;
        fc1_weights[80][25] = 16'sd-61;
        fc1_weights[80][26] = 16'sd-1;
        fc1_weights[80][27] = 16'sd-52;
        fc1_weights[80][28] = 16'sd-18;
        fc1_weights[80][29] = 16'sd-5;
        fc1_weights[80][30] = 16'sd-59;
        fc1_weights[80][31] = 16'sd-69;
        fc1_weights[80][32] = 16'sd-20;
        fc1_weights[80][33] = 16'sd28;
        fc1_weights[80][34] = 16'sd-12;
        fc1_weights[80][35] = 16'sd19;
        fc1_weights[80][36] = 16'sd-90;
        fc1_weights[80][37] = 16'sd-83;
        fc1_weights[80][38] = 16'sd-58;
        fc1_weights[80][39] = 16'sd12;
        fc1_weights[80][40] = 16'sd-131;
        fc1_weights[80][41] = 16'sd12;
        fc1_weights[80][42] = 16'sd29;
        fc1_weights[80][43] = 16'sd13;
        fc1_weights[80][44] = 16'sd12;
        fc1_weights[80][45] = 16'sd88;
        fc1_weights[80][46] = 16'sd17;
        fc1_weights[80][47] = 16'sd69;
        fc1_weights[80][48] = 16'sd-44;
        fc1_weights[80][49] = 16'sd-42;
        fc1_weights[80][50] = 16'sd0;
        fc1_weights[80][51] = 16'sd64;
        fc1_weights[80][52] = 16'sd-9;
        fc1_weights[80][53] = 16'sd-20;
        fc1_weights[80][54] = 16'sd-47;
        fc1_weights[80][55] = 16'sd0;
        fc1_weights[80][56] = 16'sd-44;
        fc1_weights[80][57] = 16'sd-42;
        fc1_weights[80][58] = 16'sd10;
        fc1_weights[80][59] = 16'sd15;
        fc1_weights[80][60] = 16'sd-66;
        fc1_weights[80][61] = 16'sd-21;
        fc1_weights[80][62] = 16'sd64;
        fc1_weights[80][63] = 16'sd-55;
        fc1_weights[80][64] = 16'sd-64;
        fc1_weights[80][65] = 16'sd41;
        fc1_weights[80][66] = 16'sd-24;
        fc1_weights[80][67] = 16'sd68;
        fc1_weights[80][68] = 16'sd79;
        fc1_weights[80][69] = 16'sd40;
        fc1_weights[80][70] = 16'sd66;
        fc1_weights[80][71] = 16'sd34;
        fc1_weights[80][72] = 16'sd-1;
        fc1_weights[80][73] = 16'sd28;
        fc1_weights[80][74] = 16'sd18;
        fc1_weights[80][75] = 16'sd26;
        fc1_weights[80][76] = 16'sd-24;
        fc1_weights[80][77] = 16'sd44;
        fc1_weights[80][78] = 16'sd-56;
        fc1_weights[80][79] = 16'sd-64;
        fc1_weights[80][80] = 16'sd-62;
        fc1_weights[80][81] = 16'sd-21;
        fc1_weights[80][82] = 16'sd-4;
        fc1_weights[80][83] = 16'sd19;
        fc1_weights[80][84] = 16'sd41;
        fc1_weights[80][85] = 16'sd41;
        fc1_weights[80][86] = 16'sd16;
        fc1_weights[80][87] = 16'sd7;
        fc1_weights[80][88] = 16'sd59;
        fc1_weights[80][89] = 16'sd-36;
        fc1_weights[80][90] = 16'sd8;
        fc1_weights[80][91] = 16'sd-66;
        fc1_weights[80][92] = 16'sd-34;
        fc1_weights[80][93] = 16'sd-33;
        fc1_weights[80][94] = 16'sd29;
        fc1_weights[80][95] = 16'sd-3;
        fc1_weights[80][96] = 16'sd100;
        fc1_weights[80][97] = 16'sd35;
        fc1_weights[80][98] = 16'sd-9;
        fc1_weights[80][99] = 16'sd-6;
        fc1_weights[80][100] = 16'sd18;
        fc1_weights[80][101] = 16'sd38;
        fc1_weights[80][102] = 16'sd44;
        fc1_weights[80][103] = 16'sd84;
        fc1_weights[80][104] = 16'sd-40;
        fc1_weights[80][105] = 16'sd-9;
        fc1_weights[80][106] = 16'sd-6;
        fc1_weights[80][107] = 16'sd19;
        fc1_weights[80][108] = 16'sd-23;
        fc1_weights[80][109] = 16'sd-21;
        fc1_weights[80][110] = 16'sd-6;
        fc1_weights[80][111] = 16'sd16;
        fc1_weights[80][112] = 16'sd28;
        fc1_weights[80][113] = 16'sd42;
        fc1_weights[80][114] = 16'sd-31;
        fc1_weights[80][115] = 16'sd5;
        fc1_weights[80][116] = 16'sd22;
        fc1_weights[80][117] = 16'sd-3;
        fc1_weights[80][118] = 16'sd-4;
        fc1_weights[80][119] = 16'sd19;
        fc1_weights[80][120] = 16'sd14;
        fc1_weights[80][121] = 16'sd5;
        fc1_weights[80][122] = 16'sd-1;
        fc1_weights[80][123] = 16'sd54;
        fc1_weights[80][124] = 16'sd38;
        fc1_weights[80][125] = 16'sd-19;
        fc1_weights[80][126] = 16'sd52;
        fc1_weights[80][127] = 16'sd-10;
        fc1_weights[80][128] = 16'sd24;
        fc1_weights[80][129] = 16'sd56;
        fc1_weights[80][130] = 16'sd-26;
        fc1_weights[80][131] = 16'sd-12;
        fc1_weights[80][132] = 16'sd-28;
        fc1_weights[80][133] = 16'sd-6;
        fc1_weights[80][134] = 16'sd-49;
        fc1_weights[80][135] = 16'sd-59;
        fc1_weights[80][136] = 16'sd-61;
        fc1_weights[80][137] = 16'sd5;
        fc1_weights[80][138] = 16'sd-32;
        fc1_weights[80][139] = 16'sd-23;
        fc1_weights[80][140] = 16'sd-1;
        fc1_weights[80][141] = 16'sd3;
        fc1_weights[80][142] = 16'sd-7;
        fc1_weights[80][143] = 16'sd-11;
        fc1_weights[80][144] = 16'sd0;
        fc1_weights[80][145] = 16'sd60;
        fc1_weights[80][146] = 16'sd39;
        fc1_weights[80][147] = 16'sd36;
        fc1_weights[80][148] = 16'sd22;
        fc1_weights[80][149] = 16'sd49;
        fc1_weights[80][150] = 16'sd-14;
        fc1_weights[80][151] = 16'sd11;
        fc1_weights[80][152] = 16'sd-46;
        fc1_weights[80][153] = 16'sd-10;
        fc1_weights[80][154] = 16'sd-21;
        fc1_weights[80][155] = 16'sd-10;
        fc1_weights[80][156] = 16'sd-2;
        fc1_weights[80][157] = 16'sd-9;
        fc1_weights[80][158] = 16'sd17;
        fc1_weights[80][159] = 16'sd51;
        fc1_weights[80][160] = 16'sd-13;
        fc1_weights[80][161] = 16'sd-8;
        fc1_weights[80][162] = 16'sd-20;
        fc1_weights[80][163] = 16'sd-16;
        fc1_weights[80][164] = 16'sd-32;
        fc1_weights[80][165] = 16'sd-25;
        fc1_weights[80][166] = 16'sd-50;
        fc1_weights[80][167] = 16'sd-36;
        fc1_weights[80][168] = 16'sd-42;
        fc1_weights[80][169] = 16'sd-7;
        fc1_weights[80][170] = 16'sd-24;
        fc1_weights[80][171] = 16'sd-5;
        fc1_weights[80][172] = 16'sd-23;
        fc1_weights[80][173] = 16'sd7;
        fc1_weights[80][174] = 16'sd27;
        fc1_weights[80][175] = 16'sd-6;
        fc1_weights[80][176] = 16'sd5;
        fc1_weights[80][177] = 16'sd10;
        fc1_weights[80][178] = 16'sd56;
        fc1_weights[80][179] = 16'sd-12;
        fc1_weights[80][180] = 16'sd37;
        fc1_weights[80][181] = 16'sd28;
        fc1_weights[80][182] = 16'sd-17;
        fc1_weights[80][183] = 16'sd-23;
        fc1_weights[80][184] = 16'sd17;
        fc1_weights[80][185] = 16'sd-56;
        fc1_weights[80][186] = 16'sd-21;
        fc1_weights[80][187] = 16'sd-19;
        fc1_weights[80][188] = 16'sd-25;
        fc1_weights[80][189] = 16'sd-51;
        fc1_weights[80][190] = 16'sd-24;
        fc1_weights[80][191] = 16'sd-69;
        fc1_weights[80][192] = 16'sd8;
        fc1_weights[80][193] = 16'sd-13;
        fc1_weights[80][194] = 16'sd-7;
        fc1_weights[80][195] = 16'sd14;
        fc1_weights[80][196] = 16'sd38;
        fc1_weights[80][197] = 16'sd-23;
        fc1_weights[80][198] = 16'sd48;
        fc1_weights[80][199] = 16'sd3;
        fc1_weights[80][200] = 16'sd29;
        fc1_weights[80][201] = 16'sd27;
        fc1_weights[80][202] = 16'sd0;
        fc1_weights[80][203] = 16'sd8;
        fc1_weights[80][204] = 16'sd-26;
        fc1_weights[80][205] = 16'sd-24;
        fc1_weights[80][206] = 16'sd22;
        fc1_weights[80][207] = 16'sd30;
        fc1_weights[81][0] = 16'sd-23;
        fc1_weights[81][1] = 16'sd36;
        fc1_weights[81][2] = 16'sd-32;
        fc1_weights[81][3] = 16'sd-45;
        fc1_weights[81][4] = 16'sd-59;
        fc1_weights[81][5] = 16'sd33;
        fc1_weights[81][6] = 16'sd3;
        fc1_weights[81][7] = 16'sd-8;
        fc1_weights[81][8] = 16'sd-60;
        fc1_weights[81][9] = 16'sd-64;
        fc1_weights[81][10] = 16'sd-11;
        fc1_weights[81][11] = 16'sd-42;
        fc1_weights[81][12] = 16'sd-82;
        fc1_weights[81][13] = 16'sd-24;
        fc1_weights[81][14] = 16'sd67;
        fc1_weights[81][15] = 16'sd58;
        fc1_weights[81][16] = 16'sd75;
        fc1_weights[81][17] = 16'sd45;
        fc1_weights[81][18] = 16'sd12;
        fc1_weights[81][19] = 16'sd-16;
        fc1_weights[81][20] = 16'sd44;
        fc1_weights[81][21] = 16'sd24;
        fc1_weights[81][22] = 16'sd52;
        fc1_weights[81][23] = 16'sd-25;
        fc1_weights[81][24] = 16'sd58;
        fc1_weights[81][25] = 16'sd31;
        fc1_weights[81][26] = 16'sd-12;
        fc1_weights[81][27] = 16'sd-38;
        fc1_weights[81][28] = 16'sd-44;
        fc1_weights[81][29] = 16'sd17;
        fc1_weights[81][30] = 16'sd35;
        fc1_weights[81][31] = 16'sd27;
        fc1_weights[81][32] = 16'sd4;
        fc1_weights[81][33] = 16'sd-53;
        fc1_weights[81][34] = 16'sd-1;
        fc1_weights[81][35] = 16'sd-27;
        fc1_weights[81][36] = 16'sd4;
        fc1_weights[81][37] = 16'sd-22;
        fc1_weights[81][38] = 16'sd48;
        fc1_weights[81][39] = 16'sd20;
        fc1_weights[81][40] = 16'sd91;
        fc1_weights[81][41] = 16'sd58;
        fc1_weights[81][42] = 16'sd8;
        fc1_weights[81][43] = 16'sd0;
        fc1_weights[81][44] = 16'sd-20;
        fc1_weights[81][45] = 16'sd-76;
        fc1_weights[81][46] = 16'sd-25;
        fc1_weights[81][47] = 16'sd-62;
        fc1_weights[81][48] = 16'sd-69;
        fc1_weights[81][49] = 16'sd20;
        fc1_weights[81][50] = 16'sd18;
        fc1_weights[81][51] = 16'sd-48;
        fc1_weights[81][52] = 16'sd-68;
        fc1_weights[81][53] = 16'sd-38;
        fc1_weights[81][54] = 16'sd-62;
        fc1_weights[81][55] = 16'sd-28;
        fc1_weights[81][56] = 16'sd16;
        fc1_weights[81][57] = 16'sd-19;
        fc1_weights[81][58] = 16'sd39;
        fc1_weights[81][59] = 16'sd-64;
        fc1_weights[81][60] = 16'sd-48;
        fc1_weights[81][61] = 16'sd-56;
        fc1_weights[81][62] = 16'sd-34;
        fc1_weights[81][63] = 16'sd67;
        fc1_weights[81][64] = 16'sd36;
        fc1_weights[81][65] = 16'sd-28;
        fc1_weights[81][66] = 16'sd47;
        fc1_weights[81][67] = 16'sd32;
        fc1_weights[81][68] = 16'sd17;
        fc1_weights[81][69] = 16'sd-17;
        fc1_weights[81][70] = 16'sd-5;
        fc1_weights[81][71] = 16'sd4;
        fc1_weights[81][72] = 16'sd23;
        fc1_weights[81][73] = 16'sd-10;
        fc1_weights[81][74] = 16'sd-24;
        fc1_weights[81][75] = 16'sd25;
        fc1_weights[81][76] = 16'sd35;
        fc1_weights[81][77] = 16'sd27;
        fc1_weights[81][78] = 16'sd-24;
        fc1_weights[81][79] = 16'sd17;
        fc1_weights[81][80] = 16'sd9;
        fc1_weights[81][81] = 16'sd-37;
        fc1_weights[81][82] = 16'sd-67;
        fc1_weights[81][83] = 16'sd-58;
        fc1_weights[81][84] = 16'sd2;
        fc1_weights[81][85] = 16'sd-42;
        fc1_weights[81][86] = 16'sd-19;
        fc1_weights[81][87] = 16'sd-9;
        fc1_weights[81][88] = 16'sd-38;
        fc1_weights[81][89] = 16'sd-8;
        fc1_weights[81][90] = 16'sd91;
        fc1_weights[81][91] = 16'sd79;
        fc1_weights[81][92] = 16'sd23;
        fc1_weights[81][93] = 16'sd136;
        fc1_weights[81][94] = 16'sd51;
        fc1_weights[81][95] = 16'sd49;
        fc1_weights[81][96] = 16'sd-30;
        fc1_weights[81][97] = 16'sd36;
        fc1_weights[81][98] = 16'sd28;
        fc1_weights[81][99] = 16'sd-2;
        fc1_weights[81][100] = 16'sd12;
        fc1_weights[81][101] = 16'sd12;
        fc1_weights[81][102] = 16'sd27;
        fc1_weights[81][103] = 16'sd11;
        fc1_weights[81][104] = 16'sd-36;
        fc1_weights[81][105] = 16'sd-38;
        fc1_weights[81][106] = 16'sd-11;
        fc1_weights[81][107] = 16'sd-26;
        fc1_weights[81][108] = 16'sd49;
        fc1_weights[81][109] = 16'sd-20;
        fc1_weights[81][110] = 16'sd40;
        fc1_weights[81][111] = 16'sd-59;
        fc1_weights[81][112] = 16'sd-4;
        fc1_weights[81][113] = 16'sd-39;
        fc1_weights[81][114] = 16'sd-73;
        fc1_weights[81][115] = 16'sd-47;
        fc1_weights[81][116] = 16'sd-35;
        fc1_weights[81][117] = 16'sd13;
        fc1_weights[81][118] = 16'sd15;
        fc1_weights[81][119] = 16'sd55;
        fc1_weights[81][120] = 16'sd47;
        fc1_weights[81][121] = 16'sd-41;
        fc1_weights[81][122] = 16'sd-33;
        fc1_weights[81][123] = 16'sd2;
        fc1_weights[81][124] = 16'sd-62;
        fc1_weights[81][125] = 16'sd-29;
        fc1_weights[81][126] = 16'sd-57;
        fc1_weights[81][127] = 16'sd-19;
        fc1_weights[81][128] = 16'sd16;
        fc1_weights[81][129] = 16'sd-23;
        fc1_weights[81][130] = 16'sd-48;
        fc1_weights[81][131] = 16'sd-23;
        fc1_weights[81][132] = 16'sd21;
        fc1_weights[81][133] = 16'sd51;
        fc1_weights[81][134] = 16'sd70;
        fc1_weights[81][135] = 16'sd68;
        fc1_weights[81][136] = 16'sd32;
        fc1_weights[81][137] = 16'sd-8;
        fc1_weights[81][138] = 16'sd-7;
        fc1_weights[81][139] = 16'sd38;
        fc1_weights[81][140] = 16'sd58;
        fc1_weights[81][141] = 16'sd38;
        fc1_weights[81][142] = 16'sd69;
        fc1_weights[81][143] = 16'sd-17;
        fc1_weights[81][144] = 16'sd0;
        fc1_weights[81][145] = 16'sd-10;
        fc1_weights[81][146] = 16'sd-34;
        fc1_weights[81][147] = 16'sd28;
        fc1_weights[81][148] = 16'sd-7;
        fc1_weights[81][149] = 16'sd-45;
        fc1_weights[81][150] = 16'sd-9;
        fc1_weights[81][151] = 16'sd-56;
        fc1_weights[81][152] = 16'sd10;
        fc1_weights[81][153] = 16'sd15;
        fc1_weights[81][154] = 16'sd-2;
        fc1_weights[81][155] = 16'sd45;
        fc1_weights[81][156] = 16'sd8;
        fc1_weights[81][157] = 16'sd27;
        fc1_weights[81][158] = 16'sd4;
        fc1_weights[81][159] = 16'sd-49;
        fc1_weights[81][160] = 16'sd-20;
        fc1_weights[81][161] = 16'sd-27;
        fc1_weights[81][162] = 16'sd-33;
        fc1_weights[81][163] = 16'sd-4;
        fc1_weights[81][164] = 16'sd-38;
        fc1_weights[81][165] = 16'sd3;
        fc1_weights[81][166] = 16'sd12;
        fc1_weights[81][167] = 16'sd23;
        fc1_weights[81][168] = 16'sd13;
        fc1_weights[81][169] = 16'sd18;
        fc1_weights[81][170] = 16'sd47;
        fc1_weights[81][171] = 16'sd-33;
        fc1_weights[81][172] = 16'sd0;
        fc1_weights[81][173] = 16'sd74;
        fc1_weights[81][174] = 16'sd-34;
        fc1_weights[81][175] = 16'sd25;
        fc1_weights[81][176] = 16'sd45;
        fc1_weights[81][177] = 16'sd7;
        fc1_weights[81][178] = 16'sd-33;
        fc1_weights[81][179] = 16'sd21;
        fc1_weights[81][180] = 16'sd6;
        fc1_weights[81][181] = 16'sd-1;
        fc1_weights[81][182] = 16'sd46;
        fc1_weights[81][183] = 16'sd56;
        fc1_weights[81][184] = 16'sd53;
        fc1_weights[81][185] = 16'sd10;
        fc1_weights[81][186] = 16'sd-26;
        fc1_weights[81][187] = 16'sd26;
        fc1_weights[81][188] = 16'sd-63;
        fc1_weights[81][189] = 16'sd-50;
        fc1_weights[81][190] = 16'sd-2;
        fc1_weights[81][191] = 16'sd9;
        fc1_weights[81][192] = 16'sd-22;
        fc1_weights[81][193] = 16'sd-18;
        fc1_weights[81][194] = 16'sd-9;
        fc1_weights[81][195] = 16'sd31;
        fc1_weights[81][196] = 16'sd9;
        fc1_weights[81][197] = 16'sd25;
        fc1_weights[81][198] = 16'sd-32;
        fc1_weights[81][199] = 16'sd-37;
        fc1_weights[81][200] = 16'sd-69;
        fc1_weights[81][201] = 16'sd-64;
        fc1_weights[81][202] = 16'sd-15;
        fc1_weights[81][203] = 16'sd74;
        fc1_weights[81][204] = 16'sd4;
        fc1_weights[81][205] = 16'sd72;
        fc1_weights[81][206] = 16'sd5;
        fc1_weights[81][207] = 16'sd28;
        fc1_weights[82][0] = 16'sd17;
        fc1_weights[82][1] = 16'sd12;
        fc1_weights[82][2] = 16'sd15;
        fc1_weights[82][3] = 16'sd-5;
        fc1_weights[82][4] = 16'sd-14;
        fc1_weights[82][5] = 16'sd13;
        fc1_weights[82][6] = 16'sd41;
        fc1_weights[82][7] = 16'sd59;
        fc1_weights[82][8] = 16'sd24;
        fc1_weights[82][9] = 16'sd15;
        fc1_weights[82][10] = 16'sd15;
        fc1_weights[82][11] = 16'sd11;
        fc1_weights[82][12] = 16'sd18;
        fc1_weights[82][13] = 16'sd-34;
        fc1_weights[82][14] = 16'sd7;
        fc1_weights[82][15] = 16'sd-29;
        fc1_weights[82][16] = 16'sd22;
        fc1_weights[82][17] = 16'sd-21;
        fc1_weights[82][18] = 16'sd-20;
        fc1_weights[82][19] = 16'sd-10;
        fc1_weights[82][20] = 16'sd-42;
        fc1_weights[82][21] = 16'sd23;
        fc1_weights[82][22] = 16'sd-21;
        fc1_weights[82][23] = 16'sd30;
        fc1_weights[82][24] = 16'sd-35;
        fc1_weights[82][25] = 16'sd-3;
        fc1_weights[82][26] = 16'sd-8;
        fc1_weights[82][27] = 16'sd-42;
        fc1_weights[82][28] = 16'sd19;
        fc1_weights[82][29] = 16'sd12;
        fc1_weights[82][30] = 16'sd-2;
        fc1_weights[82][31] = 16'sd23;
        fc1_weights[82][32] = 16'sd11;
        fc1_weights[82][33] = 16'sd85;
        fc1_weights[82][34] = 16'sd43;
        fc1_weights[82][35] = 16'sd-3;
        fc1_weights[82][36] = 16'sd34;
        fc1_weights[82][37] = 16'sd85;
        fc1_weights[82][38] = 16'sd44;
        fc1_weights[82][39] = 16'sd13;
        fc1_weights[82][40] = 16'sd13;
        fc1_weights[82][41] = 16'sd-34;
        fc1_weights[82][42] = 16'sd-8;
        fc1_weights[82][43] = 16'sd-11;
        fc1_weights[82][44] = 16'sd-47;
        fc1_weights[82][45] = 16'sd-21;
        fc1_weights[82][46] = 16'sd-47;
        fc1_weights[82][47] = 16'sd-34;
        fc1_weights[82][48] = 16'sd-7;
        fc1_weights[82][49] = 16'sd-18;
        fc1_weights[82][50] = 16'sd-24;
        fc1_weights[82][51] = 16'sd-17;
        fc1_weights[82][52] = 16'sd28;
        fc1_weights[82][53] = 16'sd8;
        fc1_weights[82][54] = 16'sd36;
        fc1_weights[82][55] = 16'sd16;
        fc1_weights[82][56] = 16'sd26;
        fc1_weights[82][57] = 16'sd-8;
        fc1_weights[82][58] = 16'sd3;
        fc1_weights[82][59] = 16'sd-5;
        fc1_weights[82][60] = 16'sd17;
        fc1_weights[82][61] = 16'sd13;
        fc1_weights[82][62] = 16'sd24;
        fc1_weights[82][63] = 16'sd16;
        fc1_weights[82][64] = 16'sd13;
        fc1_weights[82][65] = 16'sd22;
        fc1_weights[82][66] = 16'sd-13;
        fc1_weights[82][67] = 16'sd-8;
        fc1_weights[82][68] = 16'sd-51;
        fc1_weights[82][69] = 16'sd19;
        fc1_weights[82][70] = 16'sd7;
        fc1_weights[82][71] = 16'sd-20;
        fc1_weights[82][72] = 16'sd-30;
        fc1_weights[82][73] = 16'sd-22;
        fc1_weights[82][74] = 16'sd-5;
        fc1_weights[82][75] = 16'sd13;
        fc1_weights[82][76] = 16'sd8;
        fc1_weights[82][77] = 16'sd9;
        fc1_weights[82][78] = 16'sd-32;
        fc1_weights[82][79] = 16'sd-73;
        fc1_weights[82][80] = 16'sd0;
        fc1_weights[82][81] = 16'sd-16;
        fc1_weights[82][82] = 16'sd4;
        fc1_weights[82][83] = 16'sd76;
        fc1_weights[82][84] = 16'sd54;
        fc1_weights[82][85] = 16'sd45;
        fc1_weights[82][86] = 16'sd32;
        fc1_weights[82][87] = 16'sd23;
        fc1_weights[82][88] = 16'sd-7;
        fc1_weights[82][89] = 16'sd10;
        fc1_weights[82][90] = 16'sd-27;
        fc1_weights[82][91] = 16'sd-1;
        fc1_weights[82][92] = 16'sd-4;
        fc1_weights[82][93] = 16'sd10;
        fc1_weights[82][94] = 16'sd13;
        fc1_weights[82][95] = 16'sd-4;
        fc1_weights[82][96] = 16'sd14;
        fc1_weights[82][97] = 16'sd7;
        fc1_weights[82][98] = 16'sd-11;
        fc1_weights[82][99] = 16'sd17;
        fc1_weights[82][100] = 16'sd-4;
        fc1_weights[82][101] = 16'sd39;
        fc1_weights[82][102] = 16'sd-13;
        fc1_weights[82][103] = 16'sd7;
        fc1_weights[82][104] = 16'sd-36;
        fc1_weights[82][105] = 16'sd8;
        fc1_weights[82][106] = 16'sd11;
        fc1_weights[82][107] = 16'sd-17;
        fc1_weights[82][108] = 16'sd-3;
        fc1_weights[82][109] = 16'sd16;
        fc1_weights[82][110] = 16'sd-4;
        fc1_weights[82][111] = 16'sd59;
        fc1_weights[82][112] = 16'sd-27;
        fc1_weights[82][113] = 16'sd-25;
        fc1_weights[82][114] = 16'sd11;
        fc1_weights[82][115] = 16'sd41;
        fc1_weights[82][116] = 16'sd-17;
        fc1_weights[82][117] = 16'sd-50;
        fc1_weights[82][118] = 16'sd-18;
        fc1_weights[82][119] = 16'sd-39;
        fc1_weights[82][120] = 16'sd-20;
        fc1_weights[82][121] = 16'sd-19;
        fc1_weights[82][122] = 16'sd-14;
        fc1_weights[82][123] = 16'sd-52;
        fc1_weights[82][124] = 16'sd-24;
        fc1_weights[82][125] = 16'sd-26;
        fc1_weights[82][126] = 16'sd8;
        fc1_weights[82][127] = 16'sd-6;
        fc1_weights[82][128] = 16'sd-18;
        fc1_weights[82][129] = 16'sd34;
        fc1_weights[82][130] = 16'sd-5;
        fc1_weights[82][131] = 16'sd30;
        fc1_weights[82][132] = 16'sd-11;
        fc1_weights[82][133] = 16'sd-29;
        fc1_weights[82][134] = 16'sd-14;
        fc1_weights[82][135] = 16'sd-19;
        fc1_weights[82][136] = 16'sd-13;
        fc1_weights[82][137] = 16'sd-9;
        fc1_weights[82][138] = 16'sd9;
        fc1_weights[82][139] = 16'sd-24;
        fc1_weights[82][140] = 16'sd-2;
        fc1_weights[82][141] = 16'sd10;
        fc1_weights[82][142] = 16'sd1;
        fc1_weights[82][143] = 16'sd33;
        fc1_weights[82][144] = 16'sd-13;
        fc1_weights[82][145] = 16'sd-11;
        fc1_weights[82][146] = 16'sd0;
        fc1_weights[82][147] = 16'sd-26;
        fc1_weights[82][148] = 16'sd-35;
        fc1_weights[82][149] = 16'sd-23;
        fc1_weights[82][150] = 16'sd-12;
        fc1_weights[82][151] = 16'sd-37;
        fc1_weights[82][152] = 16'sd-3;
        fc1_weights[82][153] = 16'sd-34;
        fc1_weights[82][154] = 16'sd-30;
        fc1_weights[82][155] = 16'sd-39;
        fc1_weights[82][156] = 16'sd9;
        fc1_weights[82][157] = 16'sd-3;
        fc1_weights[82][158] = 16'sd11;
        fc1_weights[82][159] = 16'sd-14;
        fc1_weights[82][160] = 16'sd70;
        fc1_weights[82][161] = 16'sd-2;
        fc1_weights[82][162] = 16'sd38;
        fc1_weights[82][163] = 16'sd8;
        fc1_weights[82][164] = 16'sd12;
        fc1_weights[82][165] = 16'sd21;
        fc1_weights[82][166] = 16'sd21;
        fc1_weights[82][167] = 16'sd15;
        fc1_weights[82][168] = 16'sd31;
        fc1_weights[82][169] = 16'sd10;
        fc1_weights[82][170] = 16'sd-54;
        fc1_weights[82][171] = 16'sd-9;
        fc1_weights[82][172] = 16'sd19;
        fc1_weights[82][173] = 16'sd-17;
        fc1_weights[82][174] = 16'sd2;
        fc1_weights[82][175] = 16'sd-14;
        fc1_weights[82][176] = 16'sd-23;
        fc1_weights[82][177] = 16'sd-66;
        fc1_weights[82][178] = 16'sd-36;
        fc1_weights[82][179] = 16'sd-8;
        fc1_weights[82][180] = 16'sd-32;
        fc1_weights[82][181] = 16'sd-14;
        fc1_weights[82][182] = 16'sd12;
        fc1_weights[82][183] = 16'sd-2;
        fc1_weights[82][184] = 16'sd-9;
        fc1_weights[82][185] = 16'sd2;
        fc1_weights[82][186] = 16'sd25;
        fc1_weights[82][187] = 16'sd15;
        fc1_weights[82][188] = 16'sd18;
        fc1_weights[82][189] = 16'sd2;
        fc1_weights[82][190] = 16'sd-27;
        fc1_weights[82][191] = 16'sd20;
        fc1_weights[82][192] = 16'sd43;
        fc1_weights[82][193] = 16'sd31;
        fc1_weights[82][194] = 16'sd-3;
        fc1_weights[82][195] = 16'sd-11;
        fc1_weights[82][196] = 16'sd-13;
        fc1_weights[82][197] = 16'sd-41;
        fc1_weights[82][198] = 16'sd3;
        fc1_weights[82][199] = 16'sd-26;
        fc1_weights[82][200] = 16'sd-4;
        fc1_weights[82][201] = 16'sd-22;
        fc1_weights[82][202] = 16'sd-27;
        fc1_weights[82][203] = 16'sd-32;
        fc1_weights[82][204] = 16'sd8;
        fc1_weights[82][205] = 16'sd-28;
        fc1_weights[82][206] = 16'sd-32;
        fc1_weights[82][207] = 16'sd-18;
        fc1_weights[83][0] = 16'sd24;
        fc1_weights[83][1] = 16'sd2;
        fc1_weights[83][2] = 16'sd-27;
        fc1_weights[83][3] = 16'sd2;
        fc1_weights[83][4] = 16'sd3;
        fc1_weights[83][5] = 16'sd18;
        fc1_weights[83][6] = 16'sd21;
        fc1_weights[83][7] = 16'sd-9;
        fc1_weights[83][8] = 16'sd-16;
        fc1_weights[83][9] = 16'sd-8;
        fc1_weights[83][10] = 16'sd-21;
        fc1_weights[83][11] = 16'sd-24;
        fc1_weights[83][12] = 16'sd-39;
        fc1_weights[83][13] = 16'sd19;
        fc1_weights[83][14] = 16'sd-24;
        fc1_weights[83][15] = 16'sd43;
        fc1_weights[83][16] = 16'sd-8;
        fc1_weights[83][17] = 16'sd-21;
        fc1_weights[83][18] = 16'sd-19;
        fc1_weights[83][19] = 16'sd23;
        fc1_weights[83][20] = 16'sd2;
        fc1_weights[83][21] = 16'sd11;
        fc1_weights[83][22] = 16'sd2;
        fc1_weights[83][23] = 16'sd39;
        fc1_weights[83][24] = 16'sd14;
        fc1_weights[83][25] = 16'sd2;
        fc1_weights[83][26] = 16'sd29;
        fc1_weights[83][27] = 16'sd5;
        fc1_weights[83][28] = 16'sd-9;
        fc1_weights[83][29] = 16'sd-7;
        fc1_weights[83][30] = 16'sd-17;
        fc1_weights[83][31] = 16'sd8;
        fc1_weights[83][32] = 16'sd49;
        fc1_weights[83][33] = 16'sd-27;
        fc1_weights[83][34] = 16'sd-30;
        fc1_weights[83][35] = 16'sd10;
        fc1_weights[83][36] = 16'sd4;
        fc1_weights[83][37] = 16'sd-88;
        fc1_weights[83][38] = 16'sd20;
        fc1_weights[83][39] = 16'sd-11;
        fc1_weights[83][40] = 16'sd-20;
        fc1_weights[83][41] = 16'sd68;
        fc1_weights[83][42] = 16'sd3;
        fc1_weights[83][43] = 16'sd-14;
        fc1_weights[83][44] = 16'sd26;
        fc1_weights[83][45] = 16'sd41;
        fc1_weights[83][46] = 16'sd23;
        fc1_weights[83][47] = 16'sd7;
        fc1_weights[83][48] = 16'sd40;
        fc1_weights[83][49] = 16'sd52;
        fc1_weights[83][50] = 16'sd-1;
        fc1_weights[83][51] = 16'sd19;
        fc1_weights[83][52] = 16'sd15;
        fc1_weights[83][53] = 16'sd15;
        fc1_weights[83][54] = 16'sd15;
        fc1_weights[83][55] = 16'sd-18;
        fc1_weights[83][56] = 16'sd17;
        fc1_weights[83][57] = 16'sd20;
        fc1_weights[83][58] = 16'sd12;
        fc1_weights[83][59] = 16'sd21;
        fc1_weights[83][60] = 16'sd43;
        fc1_weights[83][61] = 16'sd2;
        fc1_weights[83][62] = 16'sd-4;
        fc1_weights[83][63] = 16'sd9;
        fc1_weights[83][64] = 16'sd37;
        fc1_weights[83][65] = 16'sd-34;
        fc1_weights[83][66] = 16'sd-25;
        fc1_weights[83][67] = 16'sd-3;
        fc1_weights[83][68] = 16'sd8;
        fc1_weights[83][69] = 16'sd-11;
        fc1_weights[83][70] = 16'sd-6;
        fc1_weights[83][71] = 16'sd6;
        fc1_weights[83][72] = 16'sd-25;
        fc1_weights[83][73] = 16'sd48;
        fc1_weights[83][74] = 16'sd31;
        fc1_weights[83][75] = 16'sd-2;
        fc1_weights[83][76] = 16'sd23;
        fc1_weights[83][77] = 16'sd4;
        fc1_weights[83][78] = 16'sd32;
        fc1_weights[83][79] = 16'sd27;
        fc1_weights[83][80] = 16'sd-12;
        fc1_weights[83][81] = 16'sd31;
        fc1_weights[83][82] = 16'sd5;
        fc1_weights[83][83] = 16'sd24;
        fc1_weights[83][84] = 16'sd-31;
        fc1_weights[83][85] = 16'sd7;
        fc1_weights[83][86] = 16'sd4;
        fc1_weights[83][87] = 16'sd17;
        fc1_weights[83][88] = 16'sd35;
        fc1_weights[83][89] = 16'sd3;
        fc1_weights[83][90] = 16'sd55;
        fc1_weights[83][91] = 16'sd21;
        fc1_weights[83][92] = 16'sd-33;
        fc1_weights[83][93] = 16'sd-45;
        fc1_weights[83][94] = 16'sd-24;
        fc1_weights[83][95] = 16'sd16;
        fc1_weights[83][96] = 16'sd-39;
        fc1_weights[83][97] = 16'sd-8;
        fc1_weights[83][98] = 16'sd-24;
        fc1_weights[83][99] = 16'sd6;
        fc1_weights[83][100] = 16'sd12;
        fc1_weights[83][101] = 16'sd-53;
        fc1_weights[83][102] = 16'sd-19;
        fc1_weights[83][103] = 16'sd-3;
        fc1_weights[83][104] = 16'sd51;
        fc1_weights[83][105] = 16'sd5;
        fc1_weights[83][106] = 16'sd26;
        fc1_weights[83][107] = 16'sd53;
        fc1_weights[83][108] = 16'sd-26;
        fc1_weights[83][109] = 16'sd44;
        fc1_weights[83][110] = 16'sd7;
        fc1_weights[83][111] = 16'sd18;
        fc1_weights[83][112] = 16'sd53;
        fc1_weights[83][113] = 16'sd38;
        fc1_weights[83][114] = 16'sd24;
        fc1_weights[83][115] = 16'sd-16;
        fc1_weights[83][116] = 16'sd6;
        fc1_weights[83][117] = 16'sd30;
        fc1_weights[83][118] = 16'sd55;
        fc1_weights[83][119] = 16'sd11;
        fc1_weights[83][120] = 16'sd3;
        fc1_weights[83][121] = 16'sd13;
        fc1_weights[83][122] = 16'sd-36;
        fc1_weights[83][123] = 16'sd60;
        fc1_weights[83][124] = 16'sd-11;
        fc1_weights[83][125] = 16'sd45;
        fc1_weights[83][126] = 16'sd18;
        fc1_weights[83][127] = 16'sd22;
        fc1_weights[83][128] = 16'sd23;
        fc1_weights[83][129] = 16'sd44;
        fc1_weights[83][130] = 16'sd43;
        fc1_weights[83][131] = 16'sd-7;
        fc1_weights[83][132] = 16'sd23;
        fc1_weights[83][133] = 16'sd27;
        fc1_weights[83][134] = 16'sd48;
        fc1_weights[83][135] = 16'sd40;
        fc1_weights[83][136] = 16'sd40;
        fc1_weights[83][137] = 16'sd30;
        fc1_weights[83][138] = 16'sd53;
        fc1_weights[83][139] = 16'sd-1;
        fc1_weights[83][140] = 16'sd-31;
        fc1_weights[83][141] = 16'sd-71;
        fc1_weights[83][142] = 16'sd-33;
        fc1_weights[83][143] = 16'sd-39;
        fc1_weights[83][144] = 16'sd-27;
        fc1_weights[83][145] = 16'sd-24;
        fc1_weights[83][146] = 16'sd12;
        fc1_weights[83][147] = 16'sd-8;
        fc1_weights[83][148] = 16'sd-10;
        fc1_weights[83][149] = 16'sd-3;
        fc1_weights[83][150] = 16'sd-8;
        fc1_weights[83][151] = 16'sd38;
        fc1_weights[83][152] = 16'sd-36;
        fc1_weights[83][153] = 16'sd-5;
        fc1_weights[83][154] = 16'sd27;
        fc1_weights[83][155] = 16'sd2;
        fc1_weights[83][156] = 16'sd37;
        fc1_weights[83][157] = 16'sd65;
        fc1_weights[83][158] = 16'sd1;
        fc1_weights[83][159] = 16'sd3;
        fc1_weights[83][160] = 16'sd-38;
        fc1_weights[83][161] = 16'sd15;
        fc1_weights[83][162] = 16'sd24;
        fc1_weights[83][163] = 16'sd19;
        fc1_weights[83][164] = 16'sd0;
        fc1_weights[83][165] = 16'sd-46;
        fc1_weights[83][166] = 16'sd-64;
        fc1_weights[83][167] = 16'sd-32;
        fc1_weights[83][168] = 16'sd-2;
        fc1_weights[83][169] = 16'sd18;
        fc1_weights[83][170] = 16'sd23;
        fc1_weights[83][171] = 16'sd-28;
        fc1_weights[83][172] = 16'sd-49;
        fc1_weights[83][173] = 16'sd-38;
        fc1_weights[83][174] = 16'sd-25;
        fc1_weights[83][175] = 16'sd-7;
        fc1_weights[83][176] = 16'sd-42;
        fc1_weights[83][177] = 16'sd-30;
        fc1_weights[83][178] = 16'sd-5;
        fc1_weights[83][179] = 16'sd3;
        fc1_weights[83][180] = 16'sd34;
        fc1_weights[83][181] = 16'sd-1;
        fc1_weights[83][182] = 16'sd-26;
        fc1_weights[83][183] = 16'sd3;
        fc1_weights[83][184] = 16'sd45;
        fc1_weights[83][185] = 16'sd22;
        fc1_weights[83][186] = 16'sd22;
        fc1_weights[83][187] = 16'sd28;
        fc1_weights[83][188] = 16'sd11;
        fc1_weights[83][189] = 16'sd66;
        fc1_weights[83][190] = 16'sd33;
        fc1_weights[83][191] = 16'sd-26;
        fc1_weights[83][192] = 16'sd-5;
        fc1_weights[83][193] = 16'sd-25;
        fc1_weights[83][194] = 16'sd-1;
        fc1_weights[83][195] = 16'sd15;
        fc1_weights[83][196] = 16'sd27;
        fc1_weights[83][197] = 16'sd12;
        fc1_weights[83][198] = 16'sd-26;
        fc1_weights[83][199] = 16'sd7;
        fc1_weights[83][200] = 16'sd-8;
        fc1_weights[83][201] = 16'sd-13;
        fc1_weights[83][202] = 16'sd-42;
        fc1_weights[83][203] = 16'sd-9;
        fc1_weights[83][204] = 16'sd-22;
        fc1_weights[83][205] = 16'sd-26;
        fc1_weights[83][206] = 16'sd-32;
        fc1_weights[83][207] = 16'sd6;
        fc1_weights[84][0] = 16'sd30;
        fc1_weights[84][1] = 16'sd12;
        fc1_weights[84][2] = 16'sd-32;
        fc1_weights[84][3] = 16'sd-5;
        fc1_weights[84][4] = 16'sd-11;
        fc1_weights[84][5] = 16'sd-15;
        fc1_weights[84][6] = 16'sd-7;
        fc1_weights[84][7] = 16'sd30;
        fc1_weights[84][8] = 16'sd22;
        fc1_weights[84][9] = 16'sd24;
        fc1_weights[84][10] = 16'sd9;
        fc1_weights[84][11] = 16'sd3;
        fc1_weights[84][12] = 16'sd6;
        fc1_weights[84][13] = 16'sd-25;
        fc1_weights[84][14] = 16'sd-15;
        fc1_weights[84][15] = 16'sd12;
        fc1_weights[84][16] = 16'sd26;
        fc1_weights[84][17] = 16'sd3;
        fc1_weights[84][18] = 16'sd-2;
        fc1_weights[84][19] = 16'sd-9;
        fc1_weights[84][20] = 16'sd-18;
        fc1_weights[84][21] = 16'sd-6;
        fc1_weights[84][22] = 16'sd-19;
        fc1_weights[84][23] = 16'sd-40;
        fc1_weights[84][24] = 16'sd-55;
        fc1_weights[84][25] = 16'sd-56;
        fc1_weights[84][26] = 16'sd-15;
        fc1_weights[84][27] = 16'sd0;
        fc1_weights[84][28] = 16'sd-21;
        fc1_weights[84][29] = 16'sd-7;
        fc1_weights[84][30] = 16'sd0;
        fc1_weights[84][31] = 16'sd0;
        fc1_weights[84][32] = 16'sd0;
        fc1_weights[84][33] = 16'sd22;
        fc1_weights[84][34] = 16'sd10;
        fc1_weights[84][35] = 16'sd-10;
        fc1_weights[84][36] = 16'sd14;
        fc1_weights[84][37] = 16'sd19;
        fc1_weights[84][38] = 16'sd7;
        fc1_weights[84][39] = 16'sd-66;
        fc1_weights[84][40] = 16'sd-17;
        fc1_weights[84][41] = 16'sd-7;
        fc1_weights[84][42] = 16'sd-22;
        fc1_weights[84][43] = 16'sd27;
        fc1_weights[84][44] = 16'sd-24;
        fc1_weights[84][45] = 16'sd-18;
        fc1_weights[84][46] = 16'sd-34;
        fc1_weights[84][47] = 16'sd-10;
        fc1_weights[84][48] = 16'sd-17;
        fc1_weights[84][49] = 16'sd-24;
        fc1_weights[84][50] = 16'sd-49;
        fc1_weights[84][51] = 16'sd-35;
        fc1_weights[84][52] = 16'sd-5;
        fc1_weights[84][53] = 16'sd-15;
        fc1_weights[84][54] = 16'sd1;
        fc1_weights[84][55] = 16'sd-27;
        fc1_weights[84][56] = 16'sd-21;
        fc1_weights[84][57] = 16'sd-26;
        fc1_weights[84][58] = 16'sd-21;
        fc1_weights[84][59] = 16'sd-25;
        fc1_weights[84][60] = 16'sd-26;
        fc1_weights[84][61] = 16'sd-7;
        fc1_weights[84][62] = 16'sd12;
        fc1_weights[84][63] = 16'sd27;
        fc1_weights[84][64] = 16'sd-2;
        fc1_weights[84][65] = 16'sd-2;
        fc1_weights[84][66] = 16'sd33;
        fc1_weights[84][67] = 16'sd4;
        fc1_weights[84][68] = 16'sd-3;
        fc1_weights[84][69] = 16'sd17;
        fc1_weights[84][70] = 16'sd-49;
        fc1_weights[84][71] = 16'sd-8;
        fc1_weights[84][72] = 16'sd-14;
        fc1_weights[84][73] = 16'sd-66;
        fc1_weights[84][74] = 16'sd-57;
        fc1_weights[84][75] = 16'sd-13;
        fc1_weights[84][76] = 16'sd-9;
        fc1_weights[84][77] = 16'sd-25;
        fc1_weights[84][78] = 16'sd19;
        fc1_weights[84][79] = 16'sd-7;
        fc1_weights[84][80] = 16'sd-33;
        fc1_weights[84][81] = 16'sd17;
        fc1_weights[84][82] = 16'sd-1;
        fc1_weights[84][83] = 16'sd-3;
        fc1_weights[84][84] = 16'sd-12;
        fc1_weights[84][85] = 16'sd-24;
        fc1_weights[84][86] = 16'sd-30;
        fc1_weights[84][87] = 16'sd-51;
        fc1_weights[84][88] = 16'sd-24;
        fc1_weights[84][89] = 16'sd52;
        fc1_weights[84][90] = 16'sd4;
        fc1_weights[84][91] = 16'sd11;
        fc1_weights[84][92] = 16'sd41;
        fc1_weights[84][93] = 16'sd37;
        fc1_weights[84][94] = 16'sd56;
        fc1_weights[84][95] = 16'sd33;
        fc1_weights[84][96] = 16'sd8;
        fc1_weights[84][97] = 16'sd3;
        fc1_weights[84][98] = 16'sd-5;
        fc1_weights[84][99] = 16'sd-3;
        fc1_weights[84][100] = 16'sd-26;
        fc1_weights[84][101] = 16'sd-13;
        fc1_weights[84][102] = 16'sd2;
        fc1_weights[84][103] = 16'sd2;
        fc1_weights[84][104] = 16'sd3;
        fc1_weights[84][105] = 16'sd-4;
        fc1_weights[84][106] = 16'sd9;
        fc1_weights[84][107] = 16'sd-11;
        fc1_weights[84][108] = 16'sd2;
        fc1_weights[84][109] = 16'sd-16;
        fc1_weights[84][110] = 16'sd-6;
        fc1_weights[84][111] = 16'sd20;
        fc1_weights[84][112] = 16'sd-15;
        fc1_weights[84][113] = 16'sd-8;
        fc1_weights[84][114] = 16'sd-11;
        fc1_weights[84][115] = 16'sd35;
        fc1_weights[84][116] = 16'sd19;
        fc1_weights[84][117] = 16'sd22;
        fc1_weights[84][118] = 16'sd16;
        fc1_weights[84][119] = 16'sd46;
        fc1_weights[84][120] = 16'sd33;
        fc1_weights[84][121] = 16'sd40;
        fc1_weights[84][122] = 16'sd25;
        fc1_weights[84][123] = 16'sd4;
        fc1_weights[84][124] = 16'sd34;
        fc1_weights[84][125] = 16'sd-15;
        fc1_weights[84][126] = 16'sd-11;
        fc1_weights[84][127] = 16'sd-23;
        fc1_weights[84][128] = 16'sd11;
        fc1_weights[84][129] = 16'sd-19;
        fc1_weights[84][130] = 16'sd-7;
        fc1_weights[84][131] = 16'sd-36;
        fc1_weights[84][132] = 16'sd-11;
        fc1_weights[84][133] = 16'sd-27;
        fc1_weights[84][134] = 16'sd-6;
        fc1_weights[84][135] = 16'sd18;
        fc1_weights[84][136] = 16'sd-4;
        fc1_weights[84][137] = 16'sd-6;
        fc1_weights[84][138] = 16'sd-17;
        fc1_weights[84][139] = 16'sd11;
        fc1_weights[84][140] = 16'sd29;
        fc1_weights[84][141] = 16'sd-11;
        fc1_weights[84][142] = 16'sd31;
        fc1_weights[84][143] = 16'sd4;
        fc1_weights[84][144] = 16'sd23;
        fc1_weights[84][145] = 16'sd24;
        fc1_weights[84][146] = 16'sd34;
        fc1_weights[84][147] = 16'sd53;
        fc1_weights[84][148] = 16'sd37;
        fc1_weights[84][149] = 16'sd42;
        fc1_weights[84][150] = 16'sd17;
        fc1_weights[84][151] = 16'sd17;
        fc1_weights[84][152] = 16'sd39;
        fc1_weights[84][153] = 16'sd-6;
        fc1_weights[84][154] = 16'sd11;
        fc1_weights[84][155] = 16'sd-8;
        fc1_weights[84][156] = 16'sd13;
        fc1_weights[84][157] = 16'sd16;
        fc1_weights[84][158] = 16'sd-12;
        fc1_weights[84][159] = 16'sd-4;
        fc1_weights[84][160] = 16'sd-34;
        fc1_weights[84][161] = 16'sd-25;
        fc1_weights[84][162] = 16'sd14;
        fc1_weights[84][163] = 16'sd1;
        fc1_weights[84][164] = 16'sd18;
        fc1_weights[84][165] = 16'sd28;
        fc1_weights[84][166] = 16'sd56;
        fc1_weights[84][167] = 16'sd13;
        fc1_weights[84][168] = 16'sd16;
        fc1_weights[84][169] = 16'sd-11;
        fc1_weights[84][170] = 16'sd1;
        fc1_weights[84][171] = 16'sd35;
        fc1_weights[84][172] = 16'sd13;
        fc1_weights[84][173] = 16'sd3;
        fc1_weights[84][174] = 16'sd8;
        fc1_weights[84][175] = 16'sd6;
        fc1_weights[84][176] = 16'sd12;
        fc1_weights[84][177] = 16'sd35;
        fc1_weights[84][178] = 16'sd27;
        fc1_weights[84][179] = 16'sd7;
        fc1_weights[84][180] = 16'sd-5;
        fc1_weights[84][181] = 16'sd5;
        fc1_weights[84][182] = 16'sd-21;
        fc1_weights[84][183] = 16'sd0;
        fc1_weights[84][184] = 16'sd-13;
        fc1_weights[84][185] = 16'sd28;
        fc1_weights[84][186] = 16'sd-19;
        fc1_weights[84][187] = 16'sd-27;
        fc1_weights[84][188] = 16'sd9;
        fc1_weights[84][189] = 16'sd5;
        fc1_weights[84][190] = 16'sd13;
        fc1_weights[84][191] = 16'sd10;
        fc1_weights[84][192] = 16'sd-3;
        fc1_weights[84][193] = 16'sd2;
        fc1_weights[84][194] = 16'sd-7;
        fc1_weights[84][195] = 16'sd-22;
        fc1_weights[84][196] = 16'sd-8;
        fc1_weights[84][197] = 16'sd-4;
        fc1_weights[84][198] = 16'sd15;
        fc1_weights[84][199] = 16'sd12;
        fc1_weights[84][200] = 16'sd-21;
        fc1_weights[84][201] = 16'sd44;
        fc1_weights[84][202] = 16'sd25;
        fc1_weights[84][203] = 16'sd22;
        fc1_weights[84][204] = 16'sd30;
        fc1_weights[84][205] = 16'sd29;
        fc1_weights[84][206] = 16'sd0;
        fc1_weights[84][207] = 16'sd-5;
        fc1_weights[85][0] = 16'sd-49;
        fc1_weights[85][1] = 16'sd-19;
        fc1_weights[85][2] = 16'sd35;
        fc1_weights[85][3] = 16'sd-2;
        fc1_weights[85][4] = 16'sd27;
        fc1_weights[85][5] = 16'sd15;
        fc1_weights[85][6] = 16'sd30;
        fc1_weights[85][7] = 16'sd28;
        fc1_weights[85][8] = 16'sd-5;
        fc1_weights[85][9] = 16'sd7;
        fc1_weights[85][10] = 16'sd-36;
        fc1_weights[85][11] = 16'sd-24;
        fc1_weights[85][12] = 16'sd-17;
        fc1_weights[85][13] = 16'sd-25;
        fc1_weights[85][14] = 16'sd-23;
        fc1_weights[85][15] = 16'sd-31;
        fc1_weights[85][16] = 16'sd-37;
        fc1_weights[85][17] = 16'sd-19;
        fc1_weights[85][18] = 16'sd-3;
        fc1_weights[85][19] = 16'sd-10;
        fc1_weights[85][20] = 16'sd19;
        fc1_weights[85][21] = 16'sd8;
        fc1_weights[85][22] = 16'sd24;
        fc1_weights[85][23] = 16'sd25;
        fc1_weights[85][24] = 16'sd16;
        fc1_weights[85][25] = 16'sd9;
        fc1_weights[85][26] = 16'sd-36;
        fc1_weights[85][27] = 16'sd0;
        fc1_weights[85][28] = 16'sd0;
        fc1_weights[85][29] = 16'sd-2;
        fc1_weights[85][30] = 16'sd-15;
        fc1_weights[85][31] = 16'sd12;
        fc1_weights[85][32] = 16'sd25;
        fc1_weights[85][33] = 16'sd-6;
        fc1_weights[85][34] = 16'sd8;
        fc1_weights[85][35] = 16'sd7;
        fc1_weights[85][36] = 16'sd-30;
        fc1_weights[85][37] = 16'sd-16;
        fc1_weights[85][38] = 16'sd-26;
        fc1_weights[85][39] = 16'sd8;
        fc1_weights[85][40] = 16'sd-33;
        fc1_weights[85][41] = 16'sd3;
        fc1_weights[85][42] = 16'sd-14;
        fc1_weights[85][43] = 16'sd-32;
        fc1_weights[85][44] = 16'sd-11;
        fc1_weights[85][45] = 16'sd6;
        fc1_weights[85][46] = 16'sd26;
        fc1_weights[85][47] = 16'sd12;
        fc1_weights[85][48] = 16'sd21;
        fc1_weights[85][49] = 16'sd52;
        fc1_weights[85][50] = 16'sd11;
        fc1_weights[85][51] = 16'sd36;
        fc1_weights[85][52] = 16'sd-20;
        fc1_weights[85][53] = 16'sd-10;
        fc1_weights[85][54] = 16'sd-5;
        fc1_weights[85][55] = 16'sd4;
        fc1_weights[85][56] = 16'sd19;
        fc1_weights[85][57] = 16'sd-11;
        fc1_weights[85][58] = 16'sd-6;
        fc1_weights[85][59] = 16'sd-14;
        fc1_weights[85][60] = 16'sd-5;
        fc1_weights[85][61] = 16'sd-3;
        fc1_weights[85][62] = 16'sd9;
        fc1_weights[85][63] = 16'sd13;
        fc1_weights[85][64] = 16'sd22;
        fc1_weights[85][65] = 16'sd-44;
        fc1_weights[85][66] = 16'sd-19;
        fc1_weights[85][67] = 16'sd9;
        fc1_weights[85][68] = 16'sd12;
        fc1_weights[85][69] = 16'sd24;
        fc1_weights[85][70] = 16'sd9;
        fc1_weights[85][71] = 16'sd42;
        fc1_weights[85][72] = 16'sd23;
        fc1_weights[85][73] = 16'sd37;
        fc1_weights[85][74] = 16'sd32;
        fc1_weights[85][75] = 16'sd8;
        fc1_weights[85][76] = 16'sd-3;
        fc1_weights[85][77] = 16'sd13;
        fc1_weights[85][78] = 16'sd-20;
        fc1_weights[85][79] = 16'sd10;
        fc1_weights[85][80] = 16'sd1;
        fc1_weights[85][81] = 16'sd13;
        fc1_weights[85][82] = 16'sd27;
        fc1_weights[85][83] = 16'sd2;
        fc1_weights[85][84] = 16'sd0;
        fc1_weights[85][85] = 16'sd24;
        fc1_weights[85][86] = 16'sd28;
        fc1_weights[85][87] = 16'sd20;
        fc1_weights[85][88] = 16'sd-3;
        fc1_weights[85][89] = 16'sd-13;
        fc1_weights[85][90] = 16'sd-21;
        fc1_weights[85][91] = 16'sd-41;
        fc1_weights[85][92] = 16'sd4;
        fc1_weights[85][93] = 16'sd-32;
        fc1_weights[85][94] = 16'sd-5;
        fc1_weights[85][95] = 16'sd-8;
        fc1_weights[85][96] = 16'sd13;
        fc1_weights[85][97] = 16'sd-24;
        fc1_weights[85][98] = 16'sd14;
        fc1_weights[85][99] = 16'sd-20;
        fc1_weights[85][100] = 16'sd23;
        fc1_weights[85][101] = 16'sd20;
        fc1_weights[85][102] = 16'sd-19;
        fc1_weights[85][103] = 16'sd0;
        fc1_weights[85][104] = 16'sd16;
        fc1_weights[85][105] = 16'sd16;
        fc1_weights[85][106] = 16'sd10;
        fc1_weights[85][107] = 16'sd2;
        fc1_weights[85][108] = 16'sd-18;
        fc1_weights[85][109] = 16'sd-3;
        fc1_weights[85][110] = 16'sd-4;
        fc1_weights[85][111] = 16'sd17;
        fc1_weights[85][112] = 16'sd-16;
        fc1_weights[85][113] = 16'sd-34;
        fc1_weights[85][114] = 16'sd-23;
        fc1_weights[85][115] = 16'sd12;
        fc1_weights[85][116] = 16'sd-6;
        fc1_weights[85][117] = 16'sd5;
        fc1_weights[85][118] = 16'sd20;
        fc1_weights[85][119] = 16'sd11;
        fc1_weights[85][120] = 16'sd19;
        fc1_weights[85][121] = 16'sd-14;
        fc1_weights[85][122] = 16'sd-27;
        fc1_weights[85][123] = 16'sd-50;
        fc1_weights[85][124] = 16'sd-2;
        fc1_weights[85][125] = 16'sd-14;
        fc1_weights[85][126] = 16'sd25;
        fc1_weights[85][127] = 16'sd-13;
        fc1_weights[85][128] = 16'sd32;
        fc1_weights[85][129] = 16'sd76;
        fc1_weights[85][130] = 16'sd18;
        fc1_weights[85][131] = 16'sd24;
        fc1_weights[85][132] = 16'sd1;
        fc1_weights[85][133] = 16'sd0;
        fc1_weights[85][134] = 16'sd10;
        fc1_weights[85][135] = 16'sd6;
        fc1_weights[85][136] = 16'sd27;
        fc1_weights[85][137] = 16'sd-10;
        fc1_weights[85][138] = 16'sd-35;
        fc1_weights[85][139] = 16'sd-38;
        fc1_weights[85][140] = 16'sd-9;
        fc1_weights[85][141] = 16'sd68;
        fc1_weights[85][142] = 16'sd14;
        fc1_weights[85][143] = 16'sd15;
        fc1_weights[85][144] = 16'sd6;
        fc1_weights[85][145] = 16'sd17;
        fc1_weights[85][146] = 16'sd19;
        fc1_weights[85][147] = 16'sd-7;
        fc1_weights[85][148] = 16'sd-25;
        fc1_weights[85][149] = 16'sd-38;
        fc1_weights[85][150] = 16'sd-19;
        fc1_weights[85][151] = 16'sd-25;
        fc1_weights[85][152] = 16'sd-5;
        fc1_weights[85][153] = 16'sd4;
        fc1_weights[85][154] = 16'sd-14;
        fc1_weights[85][155] = 16'sd-14;
        fc1_weights[85][156] = 16'sd2;
        fc1_weights[85][157] = 16'sd11;
        fc1_weights[85][158] = 16'sd14;
        fc1_weights[85][159] = 16'sd12;
        fc1_weights[85][160] = 16'sd11;
        fc1_weights[85][161] = 16'sd8;
        fc1_weights[85][162] = 16'sd-16;
        fc1_weights[85][163] = 16'sd-18;
        fc1_weights[85][164] = 16'sd-7;
        fc1_weights[85][165] = 16'sd-10;
        fc1_weights[85][166] = 16'sd7;
        fc1_weights[85][167] = 16'sd26;
        fc1_weights[85][168] = 16'sd21;
        fc1_weights[85][169] = 16'sd27;
        fc1_weights[85][170] = 16'sd24;
        fc1_weights[85][171] = 16'sd19;
        fc1_weights[85][172] = 16'sd7;
        fc1_weights[85][173] = 16'sd18;
        fc1_weights[85][174] = 16'sd26;
        fc1_weights[85][175] = 16'sd-6;
        fc1_weights[85][176] = 16'sd-12;
        fc1_weights[85][177] = 16'sd-10;
        fc1_weights[85][178] = 16'sd12;
        fc1_weights[85][179] = 16'sd3;
        fc1_weights[85][180] = 16'sd-6;
        fc1_weights[85][181] = 16'sd-1;
        fc1_weights[85][182] = 16'sd9;
        fc1_weights[85][183] = 16'sd8;
        fc1_weights[85][184] = 16'sd23;
        fc1_weights[85][185] = 16'sd-13;
        fc1_weights[85][186] = 16'sd13;
        fc1_weights[85][187] = 16'sd0;
        fc1_weights[85][188] = 16'sd-15;
        fc1_weights[85][189] = 16'sd-12;
        fc1_weights[85][190] = 16'sd-42;
        fc1_weights[85][191] = 16'sd9;
        fc1_weights[85][192] = 16'sd36;
        fc1_weights[85][193] = 16'sd8;
        fc1_weights[85][194] = 16'sd-2;
        fc1_weights[85][195] = 16'sd9;
        fc1_weights[85][196] = 16'sd19;
        fc1_weights[85][197] = 16'sd-7;
        fc1_weights[85][198] = 16'sd9;
        fc1_weights[85][199] = 16'sd8;
        fc1_weights[85][200] = 16'sd14;
        fc1_weights[85][201] = 16'sd8;
        fc1_weights[85][202] = 16'sd37;
        fc1_weights[85][203] = 16'sd-19;
        fc1_weights[85][204] = 16'sd-4;
        fc1_weights[85][205] = 16'sd0;
        fc1_weights[85][206] = 16'sd11;
        fc1_weights[85][207] = 16'sd7;
        fc1_weights[86][0] = 16'sd-9;
        fc1_weights[86][1] = 16'sd1;
        fc1_weights[86][2] = 16'sd-5;
        fc1_weights[86][3] = 16'sd-56;
        fc1_weights[86][4] = 16'sd-15;
        fc1_weights[86][5] = 16'sd-32;
        fc1_weights[86][6] = 16'sd-39;
        fc1_weights[86][7] = 16'sd-19;
        fc1_weights[86][8] = 16'sd-15;
        fc1_weights[86][9] = 16'sd-37;
        fc1_weights[86][10] = 16'sd10;
        fc1_weights[86][11] = 16'sd4;
        fc1_weights[86][12] = 16'sd9;
        fc1_weights[86][13] = 16'sd19;
        fc1_weights[86][14] = 16'sd14;
        fc1_weights[86][15] = 16'sd1;
        fc1_weights[86][16] = 16'sd29;
        fc1_weights[86][17] = 16'sd35;
        fc1_weights[86][18] = 16'sd34;
        fc1_weights[86][19] = 16'sd-2;
        fc1_weights[86][20] = 16'sd22;
        fc1_weights[86][21] = 16'sd6;
        fc1_weights[86][22] = 16'sd-22;
        fc1_weights[86][23] = 16'sd-12;
        fc1_weights[86][24] = 16'sd4;
        fc1_weights[86][25] = 16'sd12;
        fc1_weights[86][26] = 16'sd-8;
        fc1_weights[86][27] = 16'sd-5;
        fc1_weights[86][28] = 16'sd-43;
        fc1_weights[86][29] = 16'sd-11;
        fc1_weights[86][30] = 16'sd-2;
        fc1_weights[86][31] = 16'sd-7;
        fc1_weights[86][32] = 16'sd9;
        fc1_weights[86][33] = 16'sd-15;
        fc1_weights[86][34] = 16'sd23;
        fc1_weights[86][35] = 16'sd13;
        fc1_weights[86][36] = 16'sd7;
        fc1_weights[86][37] = 16'sd9;
        fc1_weights[86][38] = 16'sd31;
        fc1_weights[86][39] = 16'sd23;
        fc1_weights[86][40] = 16'sd43;
        fc1_weights[86][41] = 16'sd19;
        fc1_weights[86][42] = 16'sd42;
        fc1_weights[86][43] = 16'sd35;
        fc1_weights[86][44] = 16'sd0;
        fc1_weights[86][45] = 16'sd14;
        fc1_weights[86][46] = 16'sd6;
        fc1_weights[86][47] = 16'sd0;
        fc1_weights[86][48] = 16'sd-22;
        fc1_weights[86][49] = 16'sd-3;
        fc1_weights[86][50] = 16'sd-3;
        fc1_weights[86][51] = 16'sd8;
        fc1_weights[86][52] = 16'sd-26;
        fc1_weights[86][53] = 16'sd-13;
        fc1_weights[86][54] = 16'sd-17;
        fc1_weights[86][55] = 16'sd-3;
        fc1_weights[86][56] = 16'sd10;
        fc1_weights[86][57] = 16'sd24;
        fc1_weights[86][58] = 16'sd8;
        fc1_weights[86][59] = 16'sd-4;
        fc1_weights[86][60] = 16'sd16;
        fc1_weights[86][61] = 16'sd12;
        fc1_weights[86][62] = 16'sd1;
        fc1_weights[86][63] = 16'sd24;
        fc1_weights[86][64] = 16'sd3;
        fc1_weights[86][65] = 16'sd23;
        fc1_weights[86][66] = 16'sd27;
        fc1_weights[86][67] = 16'sd20;
        fc1_weights[86][68] = 16'sd37;
        fc1_weights[86][69] = 16'sd20;
        fc1_weights[86][70] = 16'sd6;
        fc1_weights[86][71] = 16'sd-22;
        fc1_weights[86][72] = 16'sd-4;
        fc1_weights[86][73] = 16'sd-6;
        fc1_weights[86][74] = 16'sd-1;
        fc1_weights[86][75] = 16'sd-11;
        fc1_weights[86][76] = 16'sd-13;
        fc1_weights[86][77] = 16'sd19;
        fc1_weights[86][78] = 16'sd-19;
        fc1_weights[86][79] = 16'sd-29;
        fc1_weights[86][80] = 16'sd-16;
        fc1_weights[86][81] = 16'sd-16;
        fc1_weights[86][82] = 16'sd-29;
        fc1_weights[86][83] = 16'sd-22;
        fc1_weights[86][84] = 16'sd-13;
        fc1_weights[86][85] = 16'sd-29;
        fc1_weights[86][86] = 16'sd-16;
        fc1_weights[86][87] = 16'sd0;
        fc1_weights[86][88] = 16'sd-6;
        fc1_weights[86][89] = 16'sd-9;
        fc1_weights[86][90] = 16'sd-17;
        fc1_weights[86][91] = 16'sd-5;
        fc1_weights[86][92] = 16'sd-8;
        fc1_weights[86][93] = 16'sd-2;
        fc1_weights[86][94] = 16'sd13;
        fc1_weights[86][95] = 16'sd13;
        fc1_weights[86][96] = 16'sd-1;
        fc1_weights[86][97] = 16'sd15;
        fc1_weights[86][98] = 16'sd1;
        fc1_weights[86][99] = 16'sd3;
        fc1_weights[86][100] = 16'sd-3;
        fc1_weights[86][101] = 16'sd-12;
        fc1_weights[86][102] = 16'sd-20;
        fc1_weights[86][103] = 16'sd19;
        fc1_weights[86][104] = 16'sd-18;
        fc1_weights[86][105] = 16'sd-27;
        fc1_weights[86][106] = 16'sd-20;
        fc1_weights[86][107] = 16'sd-24;
        fc1_weights[86][108] = 16'sd-10;
        fc1_weights[86][109] = 16'sd-4;
        fc1_weights[86][110] = 16'sd0;
        fc1_weights[86][111] = 16'sd-26;
        fc1_weights[86][112] = 16'sd19;
        fc1_weights[86][113] = 16'sd38;
        fc1_weights[86][114] = 16'sd23;
        fc1_weights[86][115] = 16'sd25;
        fc1_weights[86][116] = 16'sd10;
        fc1_weights[86][117] = 16'sd7;
        fc1_weights[86][118] = 16'sd7;
        fc1_weights[86][119] = 16'sd-23;
        fc1_weights[86][120] = 16'sd-6;
        fc1_weights[86][121] = 16'sd-3;
        fc1_weights[86][122] = 16'sd-3;
        fc1_weights[86][123] = 16'sd-2;
        fc1_weights[86][124] = 16'sd-2;
        fc1_weights[86][125] = 16'sd-5;
        fc1_weights[86][126] = 16'sd1;
        fc1_weights[86][127] = 16'sd4;
        fc1_weights[86][128] = 16'sd-15;
        fc1_weights[86][129] = 16'sd4;
        fc1_weights[86][130] = 16'sd-24;
        fc1_weights[86][131] = 16'sd-8;
        fc1_weights[86][132] = 16'sd-7;
        fc1_weights[86][133] = 16'sd6;
        fc1_weights[86][134] = 16'sd9;
        fc1_weights[86][135] = 16'sd-11;
        fc1_weights[86][136] = 16'sd8;
        fc1_weights[86][137] = 16'sd-24;
        fc1_weights[86][138] = 16'sd19;
        fc1_weights[86][139] = 16'sd-8;
        fc1_weights[86][140] = 16'sd8;
        fc1_weights[86][141] = 16'sd22;
        fc1_weights[86][142] = 16'sd-5;
        fc1_weights[86][143] = 16'sd10;
        fc1_weights[86][144] = 16'sd33;
        fc1_weights[86][145] = 16'sd-9;
        fc1_weights[86][146] = 16'sd14;
        fc1_weights[86][147] = 16'sd-13;
        fc1_weights[86][148] = 16'sd2;
        fc1_weights[86][149] = 16'sd2;
        fc1_weights[86][150] = 16'sd-3;
        fc1_weights[86][151] = 16'sd18;
        fc1_weights[86][152] = 16'sd-3;
        fc1_weights[86][153] = 16'sd6;
        fc1_weights[86][154] = 16'sd-2;
        fc1_weights[86][155] = 16'sd2;
        fc1_weights[86][156] = 16'sd-14;
        fc1_weights[86][157] = 16'sd-13;
        fc1_weights[86][158] = 16'sd-7;
        fc1_weights[86][159] = 16'sd8;
        fc1_weights[86][160] = 16'sd-7;
        fc1_weights[86][161] = 16'sd18;
        fc1_weights[86][162] = 16'sd16;
        fc1_weights[86][163] = 16'sd-14;
        fc1_weights[86][164] = 16'sd-25;
        fc1_weights[86][165] = 16'sd-15;
        fc1_weights[86][166] = 16'sd-5;
        fc1_weights[86][167] = 16'sd17;
        fc1_weights[86][168] = 16'sd16;
        fc1_weights[86][169] = 16'sd11;
        fc1_weights[86][170] = 16'sd29;
        fc1_weights[86][171] = 16'sd6;
        fc1_weights[86][172] = 16'sd31;
        fc1_weights[86][173] = 16'sd22;
        fc1_weights[86][174] = 16'sd0;
        fc1_weights[86][175] = 16'sd20;
        fc1_weights[86][176] = 16'sd20;
        fc1_weights[86][177] = 16'sd36;
        fc1_weights[86][178] = 16'sd10;
        fc1_weights[86][179] = 16'sd11;
        fc1_weights[86][180] = 16'sd26;
        fc1_weights[86][181] = 16'sd5;
        fc1_weights[86][182] = 16'sd9;
        fc1_weights[86][183] = 16'sd-14;
        fc1_weights[86][184] = 16'sd-3;
        fc1_weights[86][185] = 16'sd-15;
        fc1_weights[86][186] = 16'sd-11;
        fc1_weights[86][187] = 16'sd-23;
        fc1_weights[86][188] = 16'sd-12;
        fc1_weights[86][189] = 16'sd-34;
        fc1_weights[86][190] = 16'sd30;
        fc1_weights[86][191] = 16'sd16;
        fc1_weights[86][192] = 16'sd14;
        fc1_weights[86][193] = 16'sd5;
        fc1_weights[86][194] = 16'sd-7;
        fc1_weights[86][195] = 16'sd21;
        fc1_weights[86][196] = 16'sd12;
        fc1_weights[86][197] = 16'sd20;
        fc1_weights[86][198] = 16'sd8;
        fc1_weights[86][199] = 16'sd4;
        fc1_weights[86][200] = 16'sd8;
        fc1_weights[86][201] = 16'sd-15;
        fc1_weights[86][202] = 16'sd-4;
        fc1_weights[86][203] = 16'sd17;
        fc1_weights[86][204] = 16'sd18;
        fc1_weights[86][205] = 16'sd14;
        fc1_weights[86][206] = 16'sd7;
        fc1_weights[86][207] = 16'sd12;
        fc1_weights[87][0] = 16'sd61;
        fc1_weights[87][1] = 16'sd13;
        fc1_weights[87][2] = 16'sd55;
        fc1_weights[87][3] = 16'sd47;
        fc1_weights[87][4] = 16'sd38;
        fc1_weights[87][5] = 16'sd21;
        fc1_weights[87][6] = 16'sd15;
        fc1_weights[87][7] = 16'sd22;
        fc1_weights[87][8] = 16'sd0;
        fc1_weights[87][9] = 16'sd69;
        fc1_weights[87][10] = 16'sd83;
        fc1_weights[87][11] = 16'sd35;
        fc1_weights[87][12] = 16'sd-33;
        fc1_weights[87][13] = 16'sd0;
        fc1_weights[87][14] = 16'sd27;
        fc1_weights[87][15] = 16'sd-51;
        fc1_weights[87][16] = 16'sd72;
        fc1_weights[87][17] = 16'sd-59;
        fc1_weights[87][18] = 16'sd-65;
        fc1_weights[87][19] = 16'sd-23;
        fc1_weights[87][20] = 16'sd22;
        fc1_weights[87][21] = 16'sd43;
        fc1_weights[87][22] = 16'sd23;
        fc1_weights[87][23] = 16'sd-4;
        fc1_weights[87][24] = 16'sd-1;
        fc1_weights[87][25] = 16'sd2;
        fc1_weights[87][26] = 16'sd15;
        fc1_weights[87][27] = 16'sd47;
        fc1_weights[87][28] = 16'sd27;
        fc1_weights[87][29] = 16'sd-31;
        fc1_weights[87][30] = 16'sd-52;
        fc1_weights[87][31] = 16'sd-95;
        fc1_weights[87][32] = 16'sd-41;
        fc1_weights[87][33] = 16'sd61;
        fc1_weights[87][34] = 16'sd-55;
        fc1_weights[87][35] = 16'sd23;
        fc1_weights[87][36] = 16'sd48;
        fc1_weights[87][37] = 16'sd11;
        fc1_weights[87][38] = 16'sd-4;
        fc1_weights[87][39] = 16'sd113;
        fc1_weights[87][40] = 16'sd-52;
        fc1_weights[87][41] = 16'sd33;
        fc1_weights[87][42] = 16'sd-47;
        fc1_weights[87][43] = 16'sd-13;
        fc1_weights[87][44] = 16'sd26;
        fc1_weights[87][45] = 16'sd38;
        fc1_weights[87][46] = 16'sd104;
        fc1_weights[87][47] = 16'sd52;
        fc1_weights[87][48] = 16'sd25;
        fc1_weights[87][49] = 16'sd-46;
        fc1_weights[87][50] = 16'sd35;
        fc1_weights[87][51] = 16'sd68;
        fc1_weights[87][52] = 16'sd-33;
        fc1_weights[87][53] = 16'sd63;
        fc1_weights[87][54] = 16'sd-13;
        fc1_weights[87][55] = 16'sd-12;
        fc1_weights[87][56] = 16'sd-31;
        fc1_weights[87][57] = 16'sd-40;
        fc1_weights[87][58] = 16'sd70;
        fc1_weights[87][59] = 16'sd34;
        fc1_weights[87][60] = 16'sd-1;
        fc1_weights[87][61] = 16'sd56;
        fc1_weights[87][62] = 16'sd111;
        fc1_weights[87][63] = 16'sd10;
        fc1_weights[87][64] = 16'sd64;
        fc1_weights[87][65] = 16'sd125;
        fc1_weights[87][66] = 16'sd-11;
        fc1_weights[87][67] = 16'sd-41;
        fc1_weights[87][68] = 16'sd55;
        fc1_weights[87][69] = 16'sd-1;
        fc1_weights[87][70] = 16'sd60;
        fc1_weights[87][71] = 16'sd-31;
        fc1_weights[87][72] = 16'sd-10;
        fc1_weights[87][73] = 16'sd-52;
        fc1_weights[87][74] = 16'sd-32;
        fc1_weights[87][75] = 16'sd-40;
        fc1_weights[87][76] = 16'sd-28;
        fc1_weights[87][77] = 16'sd34;
        fc1_weights[87][78] = 16'sd-14;
        fc1_weights[87][79] = 16'sd-69;
        fc1_weights[87][80] = 16'sd40;
        fc1_weights[87][81] = 16'sd0;
        fc1_weights[87][82] = 16'sd3;
        fc1_weights[87][83] = 16'sd-52;
        fc1_weights[87][84] = 16'sd-15;
        fc1_weights[87][85] = 16'sd4;
        fc1_weights[87][86] = 16'sd-10;
        fc1_weights[87][87] = 16'sd-141;
        fc1_weights[87][88] = 16'sd-93;
        fc1_weights[87][89] = 16'sd-68;
        fc1_weights[87][90] = 16'sd31;
        fc1_weights[87][91] = 16'sd28;
        fc1_weights[87][92] = 16'sd5;
        fc1_weights[87][93] = 16'sd22;
        fc1_weights[87][94] = 16'sd58;
        fc1_weights[87][95] = 16'sd-54;
        fc1_weights[87][96] = 16'sd28;
        fc1_weights[87][97] = 16'sd-33;
        fc1_weights[87][98] = 16'sd-46;
        fc1_weights[87][99] = 16'sd-1;
        fc1_weights[87][100] = 16'sd-36;
        fc1_weights[87][101] = 16'sd1;
        fc1_weights[87][102] = 16'sd17;
        fc1_weights[87][103] = 16'sd-25;
        fc1_weights[87][104] = 16'sd-34;
        fc1_weights[87][105] = 16'sd18;
        fc1_weights[87][106] = 16'sd-50;
        fc1_weights[87][107] = 16'sd-9;
        fc1_weights[87][108] = 16'sd11;
        fc1_weights[87][109] = 16'sd-17;
        fc1_weights[87][110] = 16'sd-20;
        fc1_weights[87][111] = 16'sd10;
        fc1_weights[87][112] = 16'sd-37;
        fc1_weights[87][113] = 16'sd-65;
        fc1_weights[87][114] = 16'sd-9;
        fc1_weights[87][115] = 16'sd-28;
        fc1_weights[87][116] = 16'sd0;
        fc1_weights[87][117] = 16'sd-28;
        fc1_weights[87][118] = 16'sd39;
        fc1_weights[87][119] = 16'sd-21;
        fc1_weights[87][120] = 16'sd-11;
        fc1_weights[87][121] = 16'sd-37;
        fc1_weights[87][122] = 16'sd-27;
        fc1_weights[87][123] = 16'sd-138;
        fc1_weights[87][124] = 16'sd-34;
        fc1_weights[87][125] = 16'sd-41;
        fc1_weights[87][126] = 16'sd-38;
        fc1_weights[87][127] = 16'sd-66;
        fc1_weights[87][128] = 16'sd-59;
        fc1_weights[87][129] = 16'sd-45;
        fc1_weights[87][130] = 16'sd38;
        fc1_weights[87][131] = 16'sd-15;
        fc1_weights[87][132] = 16'sd-40;
        fc1_weights[87][133] = 16'sd9;
        fc1_weights[87][134] = 16'sd21;
        fc1_weights[87][135] = 16'sd50;
        fc1_weights[87][136] = 16'sd10;
        fc1_weights[87][137] = 16'sd36;
        fc1_weights[87][138] = 16'sd17;
        fc1_weights[87][139] = 16'sd69;
        fc1_weights[87][140] = 16'sd25;
        fc1_weights[87][141] = 16'sd18;
        fc1_weights[87][142] = 16'sd-52;
        fc1_weights[87][143] = 16'sd50;
        fc1_weights[87][144] = 16'sd-19;
        fc1_weights[87][145] = 16'sd70;
        fc1_weights[87][146] = 16'sd8;
        fc1_weights[87][147] = 16'sd8;
        fc1_weights[87][148] = 16'sd-16;
        fc1_weights[87][149] = 16'sd-2;
        fc1_weights[87][150] = 16'sd-51;
        fc1_weights[87][151] = 16'sd-4;
        fc1_weights[87][152] = 16'sd23;
        fc1_weights[87][153] = 16'sd-7;
        fc1_weights[87][154] = 16'sd-43;
        fc1_weights[87][155] = 16'sd-31;
        fc1_weights[87][156] = 16'sd5;
        fc1_weights[87][157] = 16'sd-11;
        fc1_weights[87][158] = 16'sd-18;
        fc1_weights[87][159] = 16'sd4;
        fc1_weights[87][160] = 16'sd61;
        fc1_weights[87][161] = 16'sd6;
        fc1_weights[87][162] = 16'sd-16;
        fc1_weights[87][163] = 16'sd-28;
        fc1_weights[87][164] = 16'sd8;
        fc1_weights[87][165] = 16'sd0;
        fc1_weights[87][166] = 16'sd11;
        fc1_weights[87][167] = 16'sd2;
        fc1_weights[87][168] = 16'sd-61;
        fc1_weights[87][169] = 16'sd-60;
        fc1_weights[87][170] = 16'sd-46;
        fc1_weights[87][171] = 16'sd-22;
        fc1_weights[87][172] = 16'sd37;
        fc1_weights[87][173] = 16'sd37;
        fc1_weights[87][174] = 16'sd-26;
        fc1_weights[87][175] = 16'sd0;
        fc1_weights[87][176] = 16'sd-10;
        fc1_weights[87][177] = 16'sd-26;
        fc1_weights[87][178] = 16'sd-5;
        fc1_weights[87][179] = 16'sd-20;
        fc1_weights[87][180] = 16'sd-89;
        fc1_weights[87][181] = 16'sd21;
        fc1_weights[87][182] = 16'sd27;
        fc1_weights[87][183] = 16'sd46;
        fc1_weights[87][184] = 16'sd42;
        fc1_weights[87][185] = 16'sd-5;
        fc1_weights[87][186] = 16'sd72;
        fc1_weights[87][187] = 16'sd30;
        fc1_weights[87][188] = 16'sd-5;
        fc1_weights[87][189] = 16'sd31;
        fc1_weights[87][190] = 16'sd-60;
        fc1_weights[87][191] = 16'sd-19;
        fc1_weights[87][192] = 16'sd6;
        fc1_weights[87][193] = 16'sd-6;
        fc1_weights[87][194] = 16'sd-44;
        fc1_weights[87][195] = 16'sd-8;
        fc1_weights[87][196] = 16'sd-19;
        fc1_weights[87][197] = 16'sd-32;
        fc1_weights[87][198] = 16'sd39;
        fc1_weights[87][199] = 16'sd13;
        fc1_weights[87][200] = 16'sd15;
        fc1_weights[87][201] = 16'sd25;
        fc1_weights[87][202] = 16'sd-8;
        fc1_weights[87][203] = 16'sd-27;
        fc1_weights[87][204] = 16'sd19;
        fc1_weights[87][205] = 16'sd15;
        fc1_weights[87][206] = 16'sd32;
        fc1_weights[87][207] = 16'sd21;
        fc1_weights[88][0] = 16'sd-2;
        fc1_weights[88][1] = 16'sd16;
        fc1_weights[88][2] = 16'sd5;
        fc1_weights[88][3] = 16'sd11;
        fc1_weights[88][4] = 16'sd13;
        fc1_weights[88][5] = 16'sd0;
        fc1_weights[88][6] = 16'sd-20;
        fc1_weights[88][7] = 16'sd7;
        fc1_weights[88][8] = 16'sd13;
        fc1_weights[88][9] = 16'sd-24;
        fc1_weights[88][10] = 16'sd31;
        fc1_weights[88][11] = 16'sd15;
        fc1_weights[88][12] = 16'sd-31;
        fc1_weights[88][13] = 16'sd-10;
        fc1_weights[88][14] = 16'sd-44;
        fc1_weights[88][15] = 16'sd-13;
        fc1_weights[88][16] = 16'sd17;
        fc1_weights[88][17] = 16'sd-11;
        fc1_weights[88][18] = 16'sd-19;
        fc1_weights[88][19] = 16'sd-29;
        fc1_weights[88][20] = 16'sd12;
        fc1_weights[88][21] = 16'sd3;
        fc1_weights[88][22] = 16'sd-30;
        fc1_weights[88][23] = 16'sd12;
        fc1_weights[88][24] = 16'sd2;
        fc1_weights[88][25] = 16'sd19;
        fc1_weights[88][26] = 16'sd-23;
        fc1_weights[88][27] = 16'sd27;
        fc1_weights[88][28] = 16'sd50;
        fc1_weights[88][29] = 16'sd35;
        fc1_weights[88][30] = 16'sd14;
        fc1_weights[88][31] = 16'sd34;
        fc1_weights[88][32] = 16'sd-4;
        fc1_weights[88][33] = 16'sd-38;
        fc1_weights[88][34] = 16'sd-2;
        fc1_weights[88][35] = 16'sd10;
        fc1_weights[88][36] = 16'sd37;
        fc1_weights[88][37] = 16'sd71;
        fc1_weights[88][38] = 16'sd14;
        fc1_weights[88][39] = 16'sd2;
        fc1_weights[88][40] = 16'sd-7;
        fc1_weights[88][41] = 16'sd-25;
        fc1_weights[88][42] = 16'sd-23;
        fc1_weights[88][43] = 16'sd-27;
        fc1_weights[88][44] = 16'sd-6;
        fc1_weights[88][45] = 16'sd-36;
        fc1_weights[88][46] = 16'sd-30;
        fc1_weights[88][47] = 16'sd4;
        fc1_weights[88][48] = 16'sd31;
        fc1_weights[88][49] = 16'sd7;
        fc1_weights[88][50] = 16'sd4;
        fc1_weights[88][51] = 16'sd-25;
        fc1_weights[88][52] = 16'sd-29;
        fc1_weights[88][53] = 16'sd25;
        fc1_weights[88][54] = 16'sd31;
        fc1_weights[88][55] = 16'sd29;
        fc1_weights[88][56] = 16'sd11;
        fc1_weights[88][57] = 16'sd48;
        fc1_weights[88][58] = 16'sd27;
        fc1_weights[88][59] = 16'sd16;
        fc1_weights[88][60] = 16'sd41;
        fc1_weights[88][61] = 16'sd51;
        fc1_weights[88][62] = 16'sd-6;
        fc1_weights[88][63] = 16'sd1;
        fc1_weights[88][64] = 16'sd13;
        fc1_weights[88][65] = 16'sd-28;
        fc1_weights[88][66] = 16'sd-40;
        fc1_weights[88][67] = 16'sd-17;
        fc1_weights[88][68] = 16'sd-11;
        fc1_weights[88][69] = 16'sd-4;
        fc1_weights[88][70] = 16'sd-28;
        fc1_weights[88][71] = 16'sd-20;
        fc1_weights[88][72] = 16'sd5;
        fc1_weights[88][73] = 16'sd16;
        fc1_weights[88][74] = 16'sd38;
        fc1_weights[88][75] = 16'sd-7;
        fc1_weights[88][76] = 16'sd16;
        fc1_weights[88][77] = 16'sd-1;
        fc1_weights[88][78] = 16'sd-13;
        fc1_weights[88][79] = 16'sd-9;
        fc1_weights[88][80] = 16'sd14;
        fc1_weights[88][81] = 16'sd25;
        fc1_weights[88][82] = 16'sd27;
        fc1_weights[88][83] = 16'sd35;
        fc1_weights[88][84] = 16'sd20;
        fc1_weights[88][85] = 16'sd0;
        fc1_weights[88][86] = 16'sd38;
        fc1_weights[88][87] = 16'sd4;
        fc1_weights[88][88] = 16'sd-18;
        fc1_weights[88][89] = 16'sd-17;
        fc1_weights[88][90] = 16'sd8;
        fc1_weights[88][91] = 16'sd-30;
        fc1_weights[88][92] = 16'sd17;
        fc1_weights[88][93] = 16'sd-32;
        fc1_weights[88][94] = 16'sd0;
        fc1_weights[88][95] = 16'sd-5;
        fc1_weights[88][96] = 16'sd-33;
        fc1_weights[88][97] = 16'sd-18;
        fc1_weights[88][98] = 16'sd-31;
        fc1_weights[88][99] = 16'sd-17;
        fc1_weights[88][100] = 16'sd11;
        fc1_weights[88][101] = 16'sd-15;
        fc1_weights[88][102] = 16'sd-7;
        fc1_weights[88][103] = 16'sd-40;
        fc1_weights[88][104] = 16'sd-17;
        fc1_weights[88][105] = 16'sd-18;
        fc1_weights[88][106] = 16'sd5;
        fc1_weights[88][107] = 16'sd-6;
        fc1_weights[88][108] = 16'sd1;
        fc1_weights[88][109] = 16'sd-33;
        fc1_weights[88][110] = 16'sd-39;
        fc1_weights[88][111] = 16'sd1;
        fc1_weights[88][112] = 16'sd1;
        fc1_weights[88][113] = 16'sd35;
        fc1_weights[88][114] = 16'sd-22;
        fc1_weights[88][115] = 16'sd-11;
        fc1_weights[88][116] = 16'sd8;
        fc1_weights[88][117] = 16'sd0;
        fc1_weights[88][118] = 16'sd-22;
        fc1_weights[88][119] = 16'sd-23;
        fc1_weights[88][120] = 16'sd-23;
        fc1_weights[88][121] = 16'sd-3;
        fc1_weights[88][122] = 16'sd-27;
        fc1_weights[88][123] = 16'sd-36;
        fc1_weights[88][124] = 16'sd-34;
        fc1_weights[88][125] = 16'sd-41;
        fc1_weights[88][126] = 16'sd-18;
        fc1_weights[88][127] = 16'sd-27;
        fc1_weights[88][128] = 16'sd-26;
        fc1_weights[88][129] = 16'sd-41;
        fc1_weights[88][130] = 16'sd-11;
        fc1_weights[88][131] = 16'sd-35;
        fc1_weights[88][132] = 16'sd-14;
        fc1_weights[88][133] = 16'sd-33;
        fc1_weights[88][134] = 16'sd-30;
        fc1_weights[88][135] = 16'sd-32;
        fc1_weights[88][136] = 16'sd-38;
        fc1_weights[88][137] = 16'sd-19;
        fc1_weights[88][138] = 16'sd26;
        fc1_weights[88][139] = 16'sd22;
        fc1_weights[88][140] = 16'sd2;
        fc1_weights[88][141] = 16'sd26;
        fc1_weights[88][142] = 16'sd12;
        fc1_weights[88][143] = 16'sd20;
        fc1_weights[88][144] = 16'sd30;
        fc1_weights[88][145] = 16'sd19;
        fc1_weights[88][146] = 16'sd1;
        fc1_weights[88][147] = 16'sd-8;
        fc1_weights[88][148] = 16'sd-13;
        fc1_weights[88][149] = 16'sd-27;
        fc1_weights[88][150] = 16'sd-28;
        fc1_weights[88][151] = 16'sd-26;
        fc1_weights[88][152] = 16'sd-12;
        fc1_weights[88][153] = 16'sd-24;
        fc1_weights[88][154] = 16'sd-16;
        fc1_weights[88][155] = 16'sd5;
        fc1_weights[88][156] = 16'sd-26;
        fc1_weights[88][157] = 16'sd-16;
        fc1_weights[88][158] = 16'sd-28;
        fc1_weights[88][159] = 16'sd-7;
        fc1_weights[88][160] = 16'sd-16;
        fc1_weights[88][161] = 16'sd-29;
        fc1_weights[88][162] = 16'sd7;
        fc1_weights[88][163] = 16'sd-29;
        fc1_weights[88][164] = 16'sd3;
        fc1_weights[88][165] = 16'sd-1;
        fc1_weights[88][166] = 16'sd-6;
        fc1_weights[88][167] = 16'sd-1;
        fc1_weights[88][168] = 16'sd5;
        fc1_weights[88][169] = 16'sd0;
        fc1_weights[88][170] = 16'sd-24;
        fc1_weights[88][171] = 16'sd8;
        fc1_weights[88][172] = 16'sd33;
        fc1_weights[88][173] = 16'sd27;
        fc1_weights[88][174] = 16'sd12;
        fc1_weights[88][175] = 16'sd-1;
        fc1_weights[88][176] = 16'sd1;
        fc1_weights[88][177] = 16'sd-4;
        fc1_weights[88][178] = 16'sd-4;
        fc1_weights[88][179] = 16'sd5;
        fc1_weights[88][180] = 16'sd0;
        fc1_weights[88][181] = 16'sd-19;
        fc1_weights[88][182] = 16'sd-18;
        fc1_weights[88][183] = 16'sd-26;
        fc1_weights[88][184] = 16'sd-31;
        fc1_weights[88][185] = 16'sd21;
        fc1_weights[88][186] = 16'sd29;
        fc1_weights[88][187] = 16'sd6;
        fc1_weights[88][188] = 16'sd-13;
        fc1_weights[88][189] = 16'sd-28;
        fc1_weights[88][190] = 16'sd29;
        fc1_weights[88][191] = 16'sd31;
        fc1_weights[88][192] = 16'sd24;
        fc1_weights[88][193] = 16'sd3;
        fc1_weights[88][194] = 16'sd18;
        fc1_weights[88][195] = 16'sd10;
        fc1_weights[88][196] = 16'sd0;
        fc1_weights[88][197] = 16'sd5;
        fc1_weights[88][198] = 16'sd-12;
        fc1_weights[88][199] = 16'sd45;
        fc1_weights[88][200] = 16'sd34;
        fc1_weights[88][201] = 16'sd27;
        fc1_weights[88][202] = 16'sd3;
        fc1_weights[88][203] = 16'sd29;
        fc1_weights[88][204] = 16'sd23;
        fc1_weights[88][205] = 16'sd-21;
        fc1_weights[88][206] = 16'sd-3;
        fc1_weights[88][207] = 16'sd-3;
        fc1_weights[89][0] = 16'sd54;
        fc1_weights[89][1] = 16'sd56;
        fc1_weights[89][2] = 16'sd12;
        fc1_weights[89][3] = 16'sd-47;
        fc1_weights[89][4] = 16'sd3;
        fc1_weights[89][5] = 16'sd35;
        fc1_weights[89][6] = 16'sd14;
        fc1_weights[89][7] = 16'sd1;
        fc1_weights[89][8] = 16'sd27;
        fc1_weights[89][9] = 16'sd-14;
        fc1_weights[89][10] = 16'sd-1;
        fc1_weights[89][11] = 16'sd-29;
        fc1_weights[89][12] = 16'sd52;
        fc1_weights[89][13] = 16'sd51;
        fc1_weights[89][14] = 16'sd60;
        fc1_weights[89][15] = 16'sd36;
        fc1_weights[89][16] = 16'sd62;
        fc1_weights[89][17] = 16'sd77;
        fc1_weights[89][18] = 16'sd17;
        fc1_weights[89][19] = 16'sd-28;
        fc1_weights[89][20] = 16'sd-35;
        fc1_weights[89][21] = 16'sd-44;
        fc1_weights[89][22] = 16'sd-9;
        fc1_weights[89][23] = 16'sd-4;
        fc1_weights[89][24] = 16'sd-67;
        fc1_weights[89][25] = 16'sd-22;
        fc1_weights[89][26] = 16'sd15;
        fc1_weights[89][27] = 16'sd4;
        fc1_weights[89][28] = 16'sd20;
        fc1_weights[89][29] = 16'sd24;
        fc1_weights[89][30] = 16'sd-33;
        fc1_weights[89][31] = 16'sd15;
        fc1_weights[89][32] = 16'sd14;
        fc1_weights[89][33] = 16'sd5;
        fc1_weights[89][34] = 16'sd30;
        fc1_weights[89][35] = 16'sd-4;
        fc1_weights[89][36] = 16'sd-50;
        fc1_weights[89][37] = 16'sd-7;
        fc1_weights[89][38] = 16'sd74;
        fc1_weights[89][39] = 16'sd16;
        fc1_weights[89][40] = 16'sd-43;
        fc1_weights[89][41] = 16'sd14;
        fc1_weights[89][42] = 16'sd40;
        fc1_weights[89][43] = 16'sd-66;
        fc1_weights[89][44] = 16'sd-15;
        fc1_weights[89][45] = 16'sd24;
        fc1_weights[89][46] = 16'sd37;
        fc1_weights[89][47] = 16'sd-9;
        fc1_weights[89][48] = 16'sd-17;
        fc1_weights[89][49] = 16'sd23;
        fc1_weights[89][50] = 16'sd19;
        fc1_weights[89][51] = 16'sd17;
        fc1_weights[89][52] = 16'sd-29;
        fc1_weights[89][53] = 16'sd-32;
        fc1_weights[89][54] = 16'sd-53;
        fc1_weights[89][55] = 16'sd-28;
        fc1_weights[89][56] = 16'sd-26;
        fc1_weights[89][57] = 16'sd-34;
        fc1_weights[89][58] = 16'sd-44;
        fc1_weights[89][59] = 16'sd6;
        fc1_weights[89][60] = 16'sd-27;
        fc1_weights[89][61] = 16'sd-48;
        fc1_weights[89][62] = 16'sd18;
        fc1_weights[89][63] = 16'sd36;
        fc1_weights[89][64] = 16'sd56;
        fc1_weights[89][65] = 16'sd-55;
        fc1_weights[89][66] = 16'sd-10;
        fc1_weights[89][67] = 16'sd-23;
        fc1_weights[89][68] = 16'sd-18;
        fc1_weights[89][69] = 16'sd29;
        fc1_weights[89][70] = 16'sd82;
        fc1_weights[89][71] = 16'sd80;
        fc1_weights[89][72] = 16'sd-4;
        fc1_weights[89][73] = 16'sd47;
        fc1_weights[89][74] = 16'sd40;
        fc1_weights[89][75] = 16'sd22;
        fc1_weights[89][76] = 16'sd-59;
        fc1_weights[89][77] = 16'sd-9;
        fc1_weights[89][78] = 16'sd-26;
        fc1_weights[89][79] = 16'sd5;
        fc1_weights[89][80] = 16'sd-55;
        fc1_weights[89][81] = 16'sd35;
        fc1_weights[89][82] = 16'sd-125;
        fc1_weights[89][83] = 16'sd-11;
        fc1_weights[89][84] = 16'sd-52;
        fc1_weights[89][85] = 16'sd2;
        fc1_weights[89][86] = 16'sd-7;
        fc1_weights[89][87] = 16'sd-5;
        fc1_weights[89][88] = 16'sd3;
        fc1_weights[89][89] = 16'sd-54;
        fc1_weights[89][90] = 16'sd23;
        fc1_weights[89][91] = 16'sd-60;
        fc1_weights[89][92] = 16'sd-12;
        fc1_weights[89][93] = 16'sd-47;
        fc1_weights[89][94] = 16'sd9;
        fc1_weights[89][95] = 16'sd65;
        fc1_weights[89][96] = 16'sd55;
        fc1_weights[89][97] = 16'sd30;
        fc1_weights[89][98] = 16'sd25;
        fc1_weights[89][99] = 16'sd-21;
        fc1_weights[89][100] = 16'sd-23;
        fc1_weights[89][101] = 16'sd-26;
        fc1_weights[89][102] = 16'sd-42;
        fc1_weights[89][103] = 16'sd-19;
        fc1_weights[89][104] = 16'sd-8;
        fc1_weights[89][105] = 16'sd-18;
        fc1_weights[89][106] = 16'sd7;
        fc1_weights[89][107] = 16'sd-24;
        fc1_weights[89][108] = 16'sd-45;
        fc1_weights[89][109] = 16'sd-5;
        fc1_weights[89][110] = 16'sd-50;
        fc1_weights[89][111] = 16'sd-58;
        fc1_weights[89][112] = 16'sd-43;
        fc1_weights[89][113] = 16'sd-65;
        fc1_weights[89][114] = 16'sd-34;
        fc1_weights[89][115] = 16'sd-31;
        fc1_weights[89][116] = 16'sd-57;
        fc1_weights[89][117] = 16'sd22;
        fc1_weights[89][118] = 16'sd-16;
        fc1_weights[89][119] = 16'sd-38;
        fc1_weights[89][120] = 16'sd10;
        fc1_weights[89][121] = 16'sd12;
        fc1_weights[89][122] = 16'sd-8;
        fc1_weights[89][123] = 16'sd-15;
        fc1_weights[89][124] = 16'sd42;
        fc1_weights[89][125] = 16'sd4;
        fc1_weights[89][126] = 16'sd16;
        fc1_weights[89][127] = 16'sd-3;
        fc1_weights[89][128] = 16'sd38;
        fc1_weights[89][129] = 16'sd31;
        fc1_weights[89][130] = 16'sd-1;
        fc1_weights[89][131] = 16'sd40;
        fc1_weights[89][132] = 16'sd-12;
        fc1_weights[89][133] = 16'sd-23;
        fc1_weights[89][134] = 16'sd-40;
        fc1_weights[89][135] = 16'sd-36;
        fc1_weights[89][136] = 16'sd-50;
        fc1_weights[89][137] = 16'sd-60;
        fc1_weights[89][138] = 16'sd-19;
        fc1_weights[89][139] = 16'sd-79;
        fc1_weights[89][140] = 16'sd-54;
        fc1_weights[89][141] = 16'sd10;
        fc1_weights[89][142] = 16'sd4;
        fc1_weights[89][143] = 16'sd-14;
        fc1_weights[89][144] = 16'sd45;
        fc1_weights[89][145] = 16'sd27;
        fc1_weights[89][146] = 16'sd3;
        fc1_weights[89][147] = 16'sd32;
        fc1_weights[89][148] = 16'sd-53;
        fc1_weights[89][149] = 16'sd-53;
        fc1_weights[89][150] = 16'sd15;
        fc1_weights[89][151] = 16'sd45;
        fc1_weights[89][152] = 16'sd-6;
        fc1_weights[89][153] = 16'sd-3;
        fc1_weights[89][154] = 16'sd47;
        fc1_weights[89][155] = 16'sd-28;
        fc1_weights[89][156] = 16'sd-21;
        fc1_weights[89][157] = 16'sd-44;
        fc1_weights[89][158] = 16'sd-27;
        fc1_weights[89][159] = 16'sd36;
        fc1_weights[89][160] = 16'sd57;
        fc1_weights[89][161] = 16'sd-15;
        fc1_weights[89][162] = 16'sd-48;
        fc1_weights[89][163] = 16'sd-24;
        fc1_weights[89][164] = 16'sd-43;
        fc1_weights[89][165] = 16'sd-35;
        fc1_weights[89][166] = 16'sd-87;
        fc1_weights[89][167] = 16'sd-59;
        fc1_weights[89][168] = 16'sd-71;
        fc1_weights[89][169] = 16'sd-14;
        fc1_weights[89][170] = 16'sd26;
        fc1_weights[89][171] = 16'sd-7;
        fc1_weights[89][172] = 16'sd-38;
        fc1_weights[89][173] = 16'sd-14;
        fc1_weights[89][174] = 16'sd-2;
        fc1_weights[89][175] = 16'sd-11;
        fc1_weights[89][176] = 16'sd-24;
        fc1_weights[89][177] = 16'sd30;
        fc1_weights[89][178] = 16'sd29;
        fc1_weights[89][179] = 16'sd-33;
        fc1_weights[89][180] = 16'sd8;
        fc1_weights[89][181] = 16'sd16;
        fc1_weights[89][182] = 16'sd-27;
        fc1_weights[89][183] = 16'sd-4;
        fc1_weights[89][184] = 16'sd10;
        fc1_weights[89][185] = 16'sd-11;
        fc1_weights[89][186] = 16'sd-16;
        fc1_weights[89][187] = 16'sd-36;
        fc1_weights[89][188] = 16'sd-17;
        fc1_weights[89][189] = 16'sd6;
        fc1_weights[89][190] = 16'sd2;
        fc1_weights[89][191] = 16'sd-82;
        fc1_weights[89][192] = 16'sd8;
        fc1_weights[89][193] = 16'sd-40;
        fc1_weights[89][194] = 16'sd29;
        fc1_weights[89][195] = 16'sd-9;
        fc1_weights[89][196] = 16'sd25;
        fc1_weights[89][197] = 16'sd-5;
        fc1_weights[89][198] = 16'sd21;
        fc1_weights[89][199] = 16'sd-9;
        fc1_weights[89][200] = 16'sd3;
        fc1_weights[89][201] = 16'sd-10;
        fc1_weights[89][202] = 16'sd-16;
        fc1_weights[89][203] = 16'sd56;
        fc1_weights[89][204] = 16'sd-78;
        fc1_weights[89][205] = 16'sd21;
        fc1_weights[89][206] = 16'sd66;
        fc1_weights[89][207] = 16'sd59;
        fc1_weights[90][0] = 16'sd26;
        fc1_weights[90][1] = 16'sd15;
        fc1_weights[90][2] = 16'sd-93;
        fc1_weights[90][3] = 16'sd19;
        fc1_weights[90][4] = 16'sd-15;
        fc1_weights[90][5] = 16'sd-13;
        fc1_weights[90][6] = 16'sd2;
        fc1_weights[90][7] = 16'sd84;
        fc1_weights[90][8] = 16'sd7;
        fc1_weights[90][9] = 16'sd-10;
        fc1_weights[90][10] = 16'sd18;
        fc1_weights[90][11] = 16'sd-18;
        fc1_weights[90][12] = 16'sd11;
        fc1_weights[90][13] = 16'sd-58;
        fc1_weights[90][14] = 16'sd-70;
        fc1_weights[90][15] = 16'sd-34;
        fc1_weights[90][16] = 16'sd-62;
        fc1_weights[90][17] = 16'sd-72;
        fc1_weights[90][18] = 16'sd39;
        fc1_weights[90][19] = 16'sd-21;
        fc1_weights[90][20] = 16'sd47;
        fc1_weights[90][21] = 16'sd-45;
        fc1_weights[90][22] = 16'sd-37;
        fc1_weights[90][23] = 16'sd-10;
        fc1_weights[90][24] = 16'sd59;
        fc1_weights[90][25] = 16'sd-32;
        fc1_weights[90][26] = 16'sd-66;
        fc1_weights[90][27] = 16'sd-28;
        fc1_weights[90][28] = 16'sd-4;
        fc1_weights[90][29] = 16'sd16;
        fc1_weights[90][30] = 16'sd18;
        fc1_weights[90][31] = 16'sd43;
        fc1_weights[90][32] = 16'sd12;
        fc1_weights[90][33] = 16'sd75;
        fc1_weights[90][34] = 16'sd-3;
        fc1_weights[90][35] = 16'sd43;
        fc1_weights[90][36] = 16'sd17;
        fc1_weights[90][37] = 16'sd88;
        fc1_weights[90][38] = 16'sd12;
        fc1_weights[90][39] = 16'sd-25;
        fc1_weights[90][40] = 16'sd6;
        fc1_weights[90][41] = 16'sd-57;
        fc1_weights[90][42] = 16'sd-20;
        fc1_weights[90][43] = 16'sd-54;
        fc1_weights[90][44] = 16'sd10;
        fc1_weights[90][45] = 16'sd-35;
        fc1_weights[90][46] = 16'sd-43;
        fc1_weights[90][47] = 16'sd-5;
        fc1_weights[90][48] = 16'sd22;
        fc1_weights[90][49] = 16'sd-15;
        fc1_weights[90][50] = 16'sd-59;
        fc1_weights[90][51] = 16'sd-25;
        fc1_weights[90][52] = 16'sd-41;
        fc1_weights[90][53] = 16'sd-75;
        fc1_weights[90][54] = 16'sd33;
        fc1_weights[90][55] = 16'sd-28;
        fc1_weights[90][56] = 16'sd-52;
        fc1_weights[90][57] = 16'sd2;
        fc1_weights[90][58] = 16'sd1;
        fc1_weights[90][59] = 16'sd16;
        fc1_weights[90][60] = 16'sd25;
        fc1_weights[90][61] = 16'sd44;
        fc1_weights[90][62] = 16'sd4;
        fc1_weights[90][63] = 16'sd12;
        fc1_weights[90][64] = 16'sd37;
        fc1_weights[90][65] = 16'sd-26;
        fc1_weights[90][66] = 16'sd-59;
        fc1_weights[90][67] = 16'sd-59;
        fc1_weights[90][68] = 16'sd-72;
        fc1_weights[90][69] = 16'sd-19;
        fc1_weights[90][70] = 16'sd-24;
        fc1_weights[90][71] = 16'sd32;
        fc1_weights[90][72] = 16'sd48;
        fc1_weights[90][73] = 16'sd-7;
        fc1_weights[90][74] = 16'sd18;
        fc1_weights[90][75] = 16'sd-36;
        fc1_weights[90][76] = 16'sd8;
        fc1_weights[90][77] = 16'sd-45;
        fc1_weights[90][78] = 16'sd36;
        fc1_weights[90][79] = 16'sd57;
        fc1_weights[90][80] = 16'sd-42;
        fc1_weights[90][81] = 16'sd18;
        fc1_weights[90][82] = 16'sd13;
        fc1_weights[90][83] = 16'sd49;
        fc1_weights[90][84] = 16'sd0;
        fc1_weights[90][85] = 16'sd-71;
        fc1_weights[90][86] = 16'sd-12;
        fc1_weights[90][87] = 16'sd35;
        fc1_weights[90][88] = 16'sd-32;
        fc1_weights[90][89] = 16'sd73;
        fc1_weights[90][90] = 16'sd12;
        fc1_weights[90][91] = 16'sd10;
        fc1_weights[90][92] = 16'sd11;
        fc1_weights[90][93] = 16'sd8;
        fc1_weights[90][94] = 16'sd-33;
        fc1_weights[90][95] = 16'sd-1;
        fc1_weights[90][96] = 16'sd17;
        fc1_weights[90][97] = 16'sd-61;
        fc1_weights[90][98] = 16'sd-5;
        fc1_weights[90][99] = 16'sd-65;
        fc1_weights[90][100] = 16'sd76;
        fc1_weights[90][101] = 16'sd1;
        fc1_weights[90][102] = 16'sd-17;
        fc1_weights[90][103] = 16'sd-29;
        fc1_weights[90][104] = 16'sd22;
        fc1_weights[90][105] = 16'sd-58;
        fc1_weights[90][106] = 16'sd-38;
        fc1_weights[90][107] = 16'sd-3;
        fc1_weights[90][108] = 16'sd8;
        fc1_weights[90][109] = 16'sd-65;
        fc1_weights[90][110] = 16'sd-36;
        fc1_weights[90][111] = 16'sd1;
        fc1_weights[90][112] = 16'sd3;
        fc1_weights[90][113] = 16'sd55;
        fc1_weights[90][114] = 16'sd30;
        fc1_weights[90][115] = 16'sd-5;
        fc1_weights[90][116] = 16'sd112;
        fc1_weights[90][117] = 16'sd67;
        fc1_weights[90][118] = 16'sd36;
        fc1_weights[90][119] = 16'sd30;
        fc1_weights[90][120] = 16'sd-29;
        fc1_weights[90][121] = 16'sd22;
        fc1_weights[90][122] = 16'sd8;
        fc1_weights[90][123] = 16'sd-43;
        fc1_weights[90][124] = 16'sd4;
        fc1_weights[90][125] = 16'sd-9;
        fc1_weights[90][126] = 16'sd15;
        fc1_weights[90][127] = 16'sd-29;
        fc1_weights[90][128] = 16'sd9;
        fc1_weights[90][129] = 16'sd-77;
        fc1_weights[90][130] = 16'sd18;
        fc1_weights[90][131] = 16'sd-33;
        fc1_weights[90][132] = 16'sd2;
        fc1_weights[90][133] = 16'sd-53;
        fc1_weights[90][134] = 16'sd-41;
        fc1_weights[90][135] = 16'sd-25;
        fc1_weights[90][136] = 16'sd-61;
        fc1_weights[90][137] = 16'sd-46;
        fc1_weights[90][138] = 16'sd4;
        fc1_weights[90][139] = 16'sd14;
        fc1_weights[90][140] = 16'sd27;
        fc1_weights[90][141] = 16'sd-92;
        fc1_weights[90][142] = 16'sd86;
        fc1_weights[90][143] = 16'sd0;
        fc1_weights[90][144] = 16'sd20;
        fc1_weights[90][145] = 16'sd57;
        fc1_weights[90][146] = 16'sd-2;
        fc1_weights[90][147] = 16'sd64;
        fc1_weights[90][148] = 16'sd46;
        fc1_weights[90][149] = 16'sd58;
        fc1_weights[90][150] = 16'sd-7;
        fc1_weights[90][151] = 16'sd20;
        fc1_weights[90][152] = 16'sd-23;
        fc1_weights[90][153] = 16'sd4;
        fc1_weights[90][154] = 16'sd-28;
        fc1_weights[90][155] = 16'sd56;
        fc1_weights[90][156] = 16'sd19;
        fc1_weights[90][157] = 16'sd-2;
        fc1_weights[90][158] = 16'sd-26;
        fc1_weights[90][159] = 16'sd63;
        fc1_weights[90][160] = 16'sd-72;
        fc1_weights[90][161] = 16'sd-69;
        fc1_weights[90][162] = 16'sd-39;
        fc1_weights[90][163] = 16'sd-3;
        fc1_weights[90][164] = 16'sd35;
        fc1_weights[90][165] = 16'sd-23;
        fc1_weights[90][166] = 16'sd75;
        fc1_weights[90][167] = 16'sd21;
        fc1_weights[90][168] = 16'sd19;
        fc1_weights[90][169] = 16'sd-14;
        fc1_weights[90][170] = 16'sd-12;
        fc1_weights[90][171] = 16'sd36;
        fc1_weights[90][172] = 16'sd21;
        fc1_weights[90][173] = 16'sd12;
        fc1_weights[90][174] = 16'sd19;
        fc1_weights[90][175] = 16'sd60;
        fc1_weights[90][176] = 16'sd30;
        fc1_weights[90][177] = 16'sd17;
        fc1_weights[90][178] = 16'sd23;
        fc1_weights[90][179] = 16'sd99;
        fc1_weights[90][180] = 16'sd40;
        fc1_weights[90][181] = 16'sd26;
        fc1_weights[90][182] = 16'sd16;
        fc1_weights[90][183] = 16'sd-16;
        fc1_weights[90][184] = 16'sd-32;
        fc1_weights[90][185] = 16'sd94;
        fc1_weights[90][186] = 16'sd-52;
        fc1_weights[90][187] = 16'sd-2;
        fc1_weights[90][188] = 16'sd2;
        fc1_weights[90][189] = 16'sd-5;
        fc1_weights[90][190] = 16'sd12;
        fc1_weights[90][191] = 16'sd54;
        fc1_weights[90][192] = 16'sd-26;
        fc1_weights[90][193] = 16'sd-9;
        fc1_weights[90][194] = 16'sd13;
        fc1_weights[90][195] = 16'sd-33;
        fc1_weights[90][196] = 16'sd-49;
        fc1_weights[90][197] = 16'sd44;
        fc1_weights[90][198] = 16'sd-9;
        fc1_weights[90][199] = 16'sd43;
        fc1_weights[90][200] = 16'sd25;
        fc1_weights[90][201] = 16'sd44;
        fc1_weights[90][202] = 16'sd25;
        fc1_weights[90][203] = 16'sd8;
        fc1_weights[90][204] = 16'sd54;
        fc1_weights[90][205] = 16'sd52;
        fc1_weights[90][206] = 16'sd6;
        fc1_weights[90][207] = 16'sd-7;
        fc1_weights[91][0] = 16'sd5;
        fc1_weights[91][1] = 16'sd-7;
        fc1_weights[91][2] = 16'sd-43;
        fc1_weights[91][3] = 16'sd5;
        fc1_weights[91][4] = 16'sd39;
        fc1_weights[91][5] = 16'sd75;
        fc1_weights[91][6] = 16'sd32;
        fc1_weights[91][7] = 16'sd19;
        fc1_weights[91][8] = 16'sd8;
        fc1_weights[91][9] = 16'sd27;
        fc1_weights[91][10] = 16'sd-25;
        fc1_weights[91][11] = 16'sd4;
        fc1_weights[91][12] = 16'sd-37;
        fc1_weights[91][13] = 16'sd-27;
        fc1_weights[91][14] = 16'sd-65;
        fc1_weights[91][15] = 16'sd-36;
        fc1_weights[91][16] = 16'sd-13;
        fc1_weights[91][17] = 16'sd9;
        fc1_weights[91][18] = 16'sd8;
        fc1_weights[91][19] = 16'sd23;
        fc1_weights[91][20] = 16'sd34;
        fc1_weights[91][21] = 16'sd-10;
        fc1_weights[91][22] = 16'sd-5;
        fc1_weights[91][23] = 16'sd52;
        fc1_weights[91][24] = 16'sd36;
        fc1_weights[91][25] = 16'sd-16;
        fc1_weights[91][26] = 16'sd-40;
        fc1_weights[91][27] = 16'sd-7;
        fc1_weights[91][28] = 16'sd-27;
        fc1_weights[91][29] = 16'sd-16;
        fc1_weights[91][30] = 16'sd17;
        fc1_weights[91][31] = 16'sd62;
        fc1_weights[91][32] = 16'sd58;
        fc1_weights[91][33] = 16'sd-40;
        fc1_weights[91][34] = 16'sd12;
        fc1_weights[91][35] = 16'sd-21;
        fc1_weights[91][36] = 16'sd39;
        fc1_weights[91][37] = 16'sd-17;
        fc1_weights[91][38] = 16'sd21;
        fc1_weights[91][39] = 16'sd20;
        fc1_weights[91][40] = 16'sd-34;
        fc1_weights[91][41] = 16'sd-16;
        fc1_weights[91][42] = 16'sd-7;
        fc1_weights[91][43] = 16'sd-17;
        fc1_weights[91][44] = 16'sd-2;
        fc1_weights[91][45] = 16'sd-11;
        fc1_weights[91][46] = 16'sd-30;
        fc1_weights[91][47] = 16'sd-48;
        fc1_weights[91][48] = 16'sd-43;
        fc1_weights[91][49] = 16'sd-18;
        fc1_weights[91][50] = 16'sd-29;
        fc1_weights[91][51] = 16'sd-6;
        fc1_weights[91][52] = 16'sd6;
        fc1_weights[91][53] = 16'sd-9;
        fc1_weights[91][54] = 16'sd18;
        fc1_weights[91][55] = 16'sd-3;
        fc1_weights[91][56] = 16'sd-15;
        fc1_weights[91][57] = 16'sd50;
        fc1_weights[91][58] = 16'sd-2;
        fc1_weights[91][59] = 16'sd35;
        fc1_weights[91][60] = 16'sd93;
        fc1_weights[91][61] = 16'sd52;
        fc1_weights[91][62] = 16'sd-30;
        fc1_weights[91][63] = 16'sd-8;
        fc1_weights[91][64] = 16'sd42;
        fc1_weights[91][65] = 16'sd37;
        fc1_weights[91][66] = 16'sd0;
        fc1_weights[91][67] = 16'sd-33;
        fc1_weights[91][68] = 16'sd-51;
        fc1_weights[91][69] = 16'sd-4;
        fc1_weights[91][70] = 16'sd-4;
        fc1_weights[91][71] = 16'sd47;
        fc1_weights[91][72] = 16'sd-13;
        fc1_weights[91][73] = 16'sd-14;
        fc1_weights[91][74] = 16'sd-17;
        fc1_weights[91][75] = 16'sd-22;
        fc1_weights[91][76] = 16'sd-3;
        fc1_weights[91][77] = 16'sd-31;
        fc1_weights[91][78] = 16'sd26;
        fc1_weights[91][79] = 16'sd40;
        fc1_weights[91][80] = 16'sd-27;
        fc1_weights[91][81] = 16'sd14;
        fc1_weights[91][82] = 16'sd-15;
        fc1_weights[91][83] = 16'sd57;
        fc1_weights[91][84] = 16'sd-28;
        fc1_weights[91][85] = 16'sd18;
        fc1_weights[91][86] = 16'sd28;
        fc1_weights[91][87] = 16'sd100;
        fc1_weights[91][88] = 16'sd10;
        fc1_weights[91][89] = 16'sd38;
        fc1_weights[91][90] = 16'sd104;
        fc1_weights[91][91] = 16'sd24;
        fc1_weights[91][92] = 16'sd-15;
        fc1_weights[91][93] = 16'sd-64;
        fc1_weights[91][94] = 16'sd-68;
        fc1_weights[91][95] = 16'sd29;
        fc1_weights[91][96] = 16'sd8;
        fc1_weights[91][97] = 16'sd3;
        fc1_weights[91][98] = 16'sd-14;
        fc1_weights[91][99] = 16'sd-19;
        fc1_weights[91][100] = 16'sd-23;
        fc1_weights[91][101] = 16'sd-17;
        fc1_weights[91][102] = 16'sd-4;
        fc1_weights[91][103] = 16'sd4;
        fc1_weights[91][104] = 16'sd27;
        fc1_weights[91][105] = 16'sd7;
        fc1_weights[91][106] = 16'sd9;
        fc1_weights[91][107] = 16'sd-2;
        fc1_weights[91][108] = 16'sd-2;
        fc1_weights[91][109] = 16'sd20;
        fc1_weights[91][110] = 16'sd-35;
        fc1_weights[91][111] = 16'sd-14;
        fc1_weights[91][112] = 16'sd18;
        fc1_weights[91][113] = 16'sd21;
        fc1_weights[91][114] = 16'sd10;
        fc1_weights[91][115] = 16'sd24;
        fc1_weights[91][116] = 16'sd45;
        fc1_weights[91][117] = 16'sd37;
        fc1_weights[91][118] = 16'sd44;
        fc1_weights[91][119] = 16'sd21;
        fc1_weights[91][120] = 16'sd18;
        fc1_weights[91][121] = 16'sd46;
        fc1_weights[91][122] = 16'sd12;
        fc1_weights[91][123] = 16'sd69;
        fc1_weights[91][124] = 16'sd6;
        fc1_weights[91][125] = 16'sd44;
        fc1_weights[91][126] = 16'sd32;
        fc1_weights[91][127] = 16'sd41;
        fc1_weights[91][128] = 16'sd25;
        fc1_weights[91][129] = 16'sd1;
        fc1_weights[91][130] = 16'sd18;
        fc1_weights[91][131] = 16'sd33;
        fc1_weights[91][132] = 16'sd3;
        fc1_weights[91][133] = 16'sd13;
        fc1_weights[91][134] = 16'sd7;
        fc1_weights[91][135] = 16'sd54;
        fc1_weights[91][136] = 16'sd-6;
        fc1_weights[91][137] = 16'sd-19;
        fc1_weights[91][138] = 16'sd-22;
        fc1_weights[91][139] = 16'sd-16;
        fc1_weights[91][140] = 16'sd-31;
        fc1_weights[91][141] = 16'sd-46;
        fc1_weights[91][142] = 16'sd10;
        fc1_weights[91][143] = 16'sd6;
        fc1_weights[91][144] = 16'sd-22;
        fc1_weights[91][145] = 16'sd-18;
        fc1_weights[91][146] = 16'sd-26;
        fc1_weights[91][147] = 16'sd3;
        fc1_weights[91][148] = 16'sd-17;
        fc1_weights[91][149] = 16'sd-17;
        fc1_weights[91][150] = 16'sd8;
        fc1_weights[91][151] = 16'sd8;
        fc1_weights[91][152] = 16'sd-41;
        fc1_weights[91][153] = 16'sd7;
        fc1_weights[91][154] = 16'sd-46;
        fc1_weights[91][155] = 16'sd29;
        fc1_weights[91][156] = 16'sd10;
        fc1_weights[91][157] = 16'sd36;
        fc1_weights[91][158] = 16'sd-39;
        fc1_weights[91][159] = 16'sd-58;
        fc1_weights[91][160] = 16'sd-57;
        fc1_weights[91][161] = 16'sd-9;
        fc1_weights[91][162] = 16'sd-4;
        fc1_weights[91][163] = 16'sd2;
        fc1_weights[91][164] = 16'sd-39;
        fc1_weights[91][165] = 16'sd-32;
        fc1_weights[91][166] = 16'sd-9;
        fc1_weights[91][167] = 16'sd-1;
        fc1_weights[91][168] = 16'sd4;
        fc1_weights[91][169] = 16'sd-5;
        fc1_weights[91][170] = 16'sd5;
        fc1_weights[91][171] = 16'sd-30;
        fc1_weights[91][172] = 16'sd-40;
        fc1_weights[91][173] = 16'sd-22;
        fc1_weights[91][174] = 16'sd-11;
        fc1_weights[91][175] = 16'sd48;
        fc1_weights[91][176] = 16'sd21;
        fc1_weights[91][177] = 16'sd-18;
        fc1_weights[91][178] = 16'sd-4;
        fc1_weights[91][179] = 16'sd10;
        fc1_weights[91][180] = 16'sd26;
        fc1_weights[91][181] = 16'sd16;
        fc1_weights[91][182] = 16'sd-18;
        fc1_weights[91][183] = 16'sd-3;
        fc1_weights[91][184] = 16'sd-17;
        fc1_weights[91][185] = 16'sd-16;
        fc1_weights[91][186] = 16'sd-19;
        fc1_weights[91][187] = 16'sd-6;
        fc1_weights[91][188] = 16'sd-31;
        fc1_weights[91][189] = 16'sd31;
        fc1_weights[91][190] = 16'sd8;
        fc1_weights[91][191] = 16'sd-9;
        fc1_weights[91][192] = 16'sd6;
        fc1_weights[91][193] = 16'sd19;
        fc1_weights[91][194] = 16'sd11;
        fc1_weights[91][195] = 16'sd1;
        fc1_weights[91][196] = 16'sd35;
        fc1_weights[91][197] = 16'sd33;
        fc1_weights[91][198] = 16'sd-23;
        fc1_weights[91][199] = 16'sd-5;
        fc1_weights[91][200] = 16'sd-23;
        fc1_weights[91][201] = 16'sd-8;
        fc1_weights[91][202] = 16'sd-42;
        fc1_weights[91][203] = 16'sd-23;
        fc1_weights[91][204] = 16'sd-10;
        fc1_weights[91][205] = 16'sd-40;
        fc1_weights[91][206] = 16'sd9;
        fc1_weights[91][207] = 16'sd-2;
        fc1_weights[92][0] = 16'sd-18;
        fc1_weights[92][1] = 16'sd17;
        fc1_weights[92][2] = 16'sd-28;
        fc1_weights[92][3] = 16'sd-80;
        fc1_weights[92][4] = 16'sd-39;
        fc1_weights[92][5] = 16'sd-5;
        fc1_weights[92][6] = 16'sd-57;
        fc1_weights[92][7] = 16'sd37;
        fc1_weights[92][8] = 16'sd-31;
        fc1_weights[92][9] = 16'sd-8;
        fc1_weights[92][10] = 16'sd75;
        fc1_weights[92][11] = 16'sd30;
        fc1_weights[92][12] = 16'sd30;
        fc1_weights[92][13] = 16'sd-25;
        fc1_weights[92][14] = 16'sd-2;
        fc1_weights[92][15] = 16'sd1;
        fc1_weights[92][16] = 16'sd-14;
        fc1_weights[92][17] = 16'sd-6;
        fc1_weights[92][18] = 16'sd-8;
        fc1_weights[92][19] = 16'sd-15;
        fc1_weights[92][20] = 16'sd42;
        fc1_weights[92][21] = 16'sd33;
        fc1_weights[92][22] = 16'sd-9;
        fc1_weights[92][23] = 16'sd-14;
        fc1_weights[92][24] = 16'sd20;
        fc1_weights[92][25] = 16'sd21;
        fc1_weights[92][26] = 16'sd-14;
        fc1_weights[92][27] = 16'sd-39;
        fc1_weights[92][28] = 16'sd-32;
        fc1_weights[92][29] = 16'sd11;
        fc1_weights[92][30] = 16'sd-18;
        fc1_weights[92][31] = 16'sd-8;
        fc1_weights[92][32] = 16'sd-16;
        fc1_weights[92][33] = 16'sd-53;
        fc1_weights[92][34] = 16'sd46;
        fc1_weights[92][35] = 16'sd58;
        fc1_weights[92][36] = 16'sd16;
        fc1_weights[92][37] = 16'sd24;
        fc1_weights[92][38] = 16'sd37;
        fc1_weights[92][39] = 16'sd0;
        fc1_weights[92][40] = 16'sd35;
        fc1_weights[92][41] = 16'sd-8;
        fc1_weights[92][42] = 16'sd-19;
        fc1_weights[92][43] = 16'sd19;
        fc1_weights[92][44] = 16'sd0;
        fc1_weights[92][45] = 16'sd32;
        fc1_weights[92][46] = 16'sd-9;
        fc1_weights[92][47] = 16'sd12;
        fc1_weights[92][48] = 16'sd6;
        fc1_weights[92][49] = 16'sd24;
        fc1_weights[92][50] = 16'sd28;
        fc1_weights[92][51] = 16'sd-11;
        fc1_weights[92][52] = 16'sd-39;
        fc1_weights[92][53] = 16'sd-49;
        fc1_weights[92][54] = 16'sd-31;
        fc1_weights[92][55] = 16'sd19;
        fc1_weights[92][56] = 16'sd17;
        fc1_weights[92][57] = 16'sd53;
        fc1_weights[92][58] = 16'sd-8;
        fc1_weights[92][59] = 16'sd-29;
        fc1_weights[92][60] = 16'sd38;
        fc1_weights[92][61] = 16'sd44;
        fc1_weights[92][62] = 16'sd-11;
        fc1_weights[92][63] = 16'sd-6;
        fc1_weights[92][64] = 16'sd79;
        fc1_weights[92][65] = 16'sd-65;
        fc1_weights[92][66] = 16'sd-13;
        fc1_weights[92][67] = 16'sd-48;
        fc1_weights[92][68] = 16'sd-74;
        fc1_weights[92][69] = 16'sd-12;
        fc1_weights[92][70] = 16'sd17;
        fc1_weights[92][71] = 16'sd9;
        fc1_weights[92][72] = 16'sd19;
        fc1_weights[92][73] = 16'sd-7;
        fc1_weights[92][74] = 16'sd42;
        fc1_weights[92][75] = 16'sd-57;
        fc1_weights[92][76] = 16'sd-32;
        fc1_weights[92][77] = 16'sd33;
        fc1_weights[92][78] = 16'sd-64;
        fc1_weights[92][79] = 16'sd-46;
        fc1_weights[92][80] = 16'sd-25;
        fc1_weights[92][81] = 16'sd-26;
        fc1_weights[92][82] = 16'sd-9;
        fc1_weights[92][83] = 16'sd8;
        fc1_weights[92][84] = 16'sd10;
        fc1_weights[92][85] = 16'sd-15;
        fc1_weights[92][86] = 16'sd-23;
        fc1_weights[92][87] = 16'sd56;
        fc1_weights[92][88] = 16'sd36;
        fc1_weights[92][89] = 16'sd-51;
        fc1_weights[92][90] = 16'sd14;
        fc1_weights[92][91] = 16'sd-2;
        fc1_weights[92][92] = 16'sd-21;
        fc1_weights[92][93] = 16'sd5;
        fc1_weights[92][94] = 16'sd-24;
        fc1_weights[92][95] = 16'sd17;
        fc1_weights[92][96] = 16'sd-30;
        fc1_weights[92][97] = 16'sd-4;
        fc1_weights[92][98] = 16'sd-2;
        fc1_weights[92][99] = 16'sd-40;
        fc1_weights[92][100] = 16'sd21;
        fc1_weights[92][101] = 16'sd-21;
        fc1_weights[92][102] = 16'sd-50;
        fc1_weights[92][103] = 16'sd-28;
        fc1_weights[92][104] = 16'sd-12;
        fc1_weights[92][105] = 16'sd-51;
        fc1_weights[92][106] = 16'sd-25;
        fc1_weights[92][107] = 16'sd-32;
        fc1_weights[92][108] = 16'sd-28;
        fc1_weights[92][109] = 16'sd-63;
        fc1_weights[92][110] = 16'sd-20;
        fc1_weights[92][111] = 16'sd20;
        fc1_weights[92][112] = 16'sd7;
        fc1_weights[92][113] = 16'sd-1;
        fc1_weights[92][114] = 16'sd56;
        fc1_weights[92][115] = 16'sd57;
        fc1_weights[92][116] = 16'sd25;
        fc1_weights[92][117] = 16'sd54;
        fc1_weights[92][118] = 16'sd60;
        fc1_weights[92][119] = 16'sd-32;
        fc1_weights[92][120] = 16'sd19;
        fc1_weights[92][121] = 16'sd32;
        fc1_weights[92][122] = 16'sd-50;
        fc1_weights[92][123] = 16'sd-28;
        fc1_weights[92][124] = 16'sd-34;
        fc1_weights[92][125] = 16'sd-28;
        fc1_weights[92][126] = 16'sd2;
        fc1_weights[92][127] = 16'sd14;
        fc1_weights[92][128] = 16'sd-48;
        fc1_weights[92][129] = 16'sd-20;
        fc1_weights[92][130] = 16'sd-15;
        fc1_weights[92][131] = 16'sd-8;
        fc1_weights[92][132] = 16'sd23;
        fc1_weights[92][133] = 16'sd-37;
        fc1_weights[92][134] = 16'sd-16;
        fc1_weights[92][135] = 16'sd-8;
        fc1_weights[92][136] = 16'sd28;
        fc1_weights[92][137] = 16'sd-32;
        fc1_weights[92][138] = 16'sd101;
        fc1_weights[92][139] = 16'sd-68;
        fc1_weights[92][140] = 16'sd-55;
        fc1_weights[92][141] = 16'sd7;
        fc1_weights[92][142] = 16'sd-21;
        fc1_weights[92][143] = 16'sd29;
        fc1_weights[92][144] = 16'sd24;
        fc1_weights[92][145] = 16'sd46;
        fc1_weights[92][146] = 16'sd4;
        fc1_weights[92][147] = 16'sd11;
        fc1_weights[92][148] = 16'sd-23;
        fc1_weights[92][149] = 16'sd7;
        fc1_weights[92][150] = 16'sd-8;
        fc1_weights[92][151] = 16'sd59;
        fc1_weights[92][152] = 16'sd-6;
        fc1_weights[92][153] = 16'sd-30;
        fc1_weights[92][154] = 16'sd-5;
        fc1_weights[92][155] = 16'sd11;
        fc1_weights[92][156] = 16'sd-49;
        fc1_weights[92][157] = 16'sd-43;
        fc1_weights[92][158] = 16'sd-31;
        fc1_weights[92][159] = 16'sd12;
        fc1_weights[92][160] = 16'sd-24;
        fc1_weights[92][161] = 16'sd18;
        fc1_weights[92][162] = 16'sd18;
        fc1_weights[92][163] = 16'sd-51;
        fc1_weights[92][164] = 16'sd-27;
        fc1_weights[92][165] = 16'sd-68;
        fc1_weights[92][166] = 16'sd0;
        fc1_weights[92][167] = 16'sd-9;
        fc1_weights[92][168] = 16'sd-20;
        fc1_weights[92][169] = 16'sd-19;
        fc1_weights[92][170] = 16'sd17;
        fc1_weights[92][171] = 16'sd-35;
        fc1_weights[92][172] = 16'sd40;
        fc1_weights[92][173] = 16'sd-3;
        fc1_weights[92][174] = 16'sd-11;
        fc1_weights[92][175] = 16'sd-29;
        fc1_weights[92][176] = 16'sd16;
        fc1_weights[92][177] = 16'sd36;
        fc1_weights[92][178] = 16'sd17;
        fc1_weights[92][179] = 16'sd67;
        fc1_weights[92][180] = 16'sd9;
        fc1_weights[92][181] = 16'sd25;
        fc1_weights[92][182] = 16'sd3;
        fc1_weights[92][183] = 16'sd-34;
        fc1_weights[92][184] = 16'sd16;
        fc1_weights[92][185] = 16'sd60;
        fc1_weights[92][186] = 16'sd3;
        fc1_weights[92][187] = 16'sd-34;
        fc1_weights[92][188] = 16'sd10;
        fc1_weights[92][189] = 16'sd-79;
        fc1_weights[92][190] = 16'sd13;
        fc1_weights[92][191] = 16'sd44;
        fc1_weights[92][192] = 16'sd33;
        fc1_weights[92][193] = 16'sd30;
        fc1_weights[92][194] = 16'sd-22;
        fc1_weights[92][195] = 16'sd30;
        fc1_weights[92][196] = 16'sd16;
        fc1_weights[92][197] = 16'sd47;
        fc1_weights[92][198] = 16'sd-25;
        fc1_weights[92][199] = 16'sd0;
        fc1_weights[92][200] = 16'sd55;
        fc1_weights[92][201] = 16'sd-10;
        fc1_weights[92][202] = 16'sd-11;
        fc1_weights[92][203] = 16'sd-19;
        fc1_weights[92][204] = 16'sd36;
        fc1_weights[92][205] = 16'sd26;
        fc1_weights[92][206] = 16'sd26;
        fc1_weights[92][207] = 16'sd47;
        fc1_weights[93][0] = 16'sd-31;
        fc1_weights[93][1] = 16'sd-33;
        fc1_weights[93][2] = 16'sd2;
        fc1_weights[93][3] = 16'sd5;
        fc1_weights[93][4] = 16'sd-21;
        fc1_weights[93][5] = 16'sd-55;
        fc1_weights[93][6] = 16'sd-22;
        fc1_weights[93][7] = 16'sd-84;
        fc1_weights[93][8] = 16'sd18;
        fc1_weights[93][9] = 16'sd45;
        fc1_weights[93][10] = 16'sd-2;
        fc1_weights[93][11] = 16'sd58;
        fc1_weights[93][12] = 16'sd45;
        fc1_weights[93][13] = 16'sd88;
        fc1_weights[93][14] = 16'sd-26;
        fc1_weights[93][15] = 16'sd-116;
        fc1_weights[93][16] = 16'sd-31;
        fc1_weights[93][17] = 16'sd-22;
        fc1_weights[93][18] = 16'sd-44;
        fc1_weights[93][19] = 16'sd-53;
        fc1_weights[93][20] = 16'sd-23;
        fc1_weights[93][21] = 16'sd-46;
        fc1_weights[93][22] = 16'sd2;
        fc1_weights[93][23] = 16'sd10;
        fc1_weights[93][24] = 16'sd-36;
        fc1_weights[93][25] = 16'sd-62;
        fc1_weights[93][26] = 16'sd91;
        fc1_weights[93][27] = 16'sd-34;
        fc1_weights[93][28] = 16'sd16;
        fc1_weights[93][29] = 16'sd-23;
        fc1_weights[93][30] = 16'sd-38;
        fc1_weights[93][31] = 16'sd-32;
        fc1_weights[93][32] = 16'sd11;
        fc1_weights[93][33] = 16'sd22;
        fc1_weights[93][34] = 16'sd-52;
        fc1_weights[93][35] = 16'sd-5;
        fc1_weights[93][36] = 16'sd4;
        fc1_weights[93][37] = 16'sd-97;
        fc1_weights[93][38] = 16'sd-7;
        fc1_weights[93][39] = 16'sd54;
        fc1_weights[93][40] = 16'sd-143;
        fc1_weights[93][41] = 16'sd-21;
        fc1_weights[93][42] = 16'sd3;
        fc1_weights[93][43] = 16'sd-19;
        fc1_weights[93][44] = 16'sd-32;
        fc1_weights[93][45] = 16'sd19;
        fc1_weights[93][46] = 16'sd17;
        fc1_weights[93][47] = 16'sd-1;
        fc1_weights[93][48] = 16'sd-56;
        fc1_weights[93][49] = 16'sd-23;
        fc1_weights[93][50] = 16'sd88;
        fc1_weights[93][51] = 16'sd90;
        fc1_weights[93][52] = 16'sd34;
        fc1_weights[93][53] = 16'sd-44;
        fc1_weights[93][54] = 16'sd-39;
        fc1_weights[93][55] = 16'sd-10;
        fc1_weights[93][56] = 16'sd-36;
        fc1_weights[93][57] = 16'sd-67;
        fc1_weights[93][58] = 16'sd25;
        fc1_weights[93][59] = 16'sd35;
        fc1_weights[93][60] = 16'sd-51;
        fc1_weights[93][61] = 16'sd-17;
        fc1_weights[93][62] = 16'sd-5;
        fc1_weights[93][63] = 16'sd1;
        fc1_weights[93][64] = 16'sd-29;
        fc1_weights[93][65] = 16'sd75;
        fc1_weights[93][66] = 16'sd-30;
        fc1_weights[93][67] = 16'sd55;
        fc1_weights[93][68] = 16'sd58;
        fc1_weights[93][69] = 16'sd0;
        fc1_weights[93][70] = 16'sd-44;
        fc1_weights[93][71] = 16'sd-22;
        fc1_weights[93][72] = 16'sd-85;
        fc1_weights[93][73] = 16'sd46;
        fc1_weights[93][74] = 16'sd-39;
        fc1_weights[93][75] = 16'sd59;
        fc1_weights[93][76] = 16'sd-4;
        fc1_weights[93][77] = 16'sd29;
        fc1_weights[93][78] = 16'sd-22;
        fc1_weights[93][79] = 16'sd-50;
        fc1_weights[93][80] = 16'sd-35;
        fc1_weights[93][81] = 16'sd-3;
        fc1_weights[93][82] = 16'sd-15;
        fc1_weights[93][83] = 16'sd-15;
        fc1_weights[93][84] = 16'sd23;
        fc1_weights[93][85] = 16'sd9;
        fc1_weights[93][86] = 16'sd53;
        fc1_weights[93][87] = 16'sd-19;
        fc1_weights[93][88] = 16'sd35;
        fc1_weights[93][89] = 16'sd-1;
        fc1_weights[93][90] = 16'sd-72;
        fc1_weights[93][91] = 16'sd-37;
        fc1_weights[93][92] = 16'sd-10;
        fc1_weights[93][93] = 16'sd46;
        fc1_weights[93][94] = 16'sd66;
        fc1_weights[93][95] = 16'sd4;
        fc1_weights[93][96] = 16'sd-28;
        fc1_weights[93][97] = 16'sd-20;
        fc1_weights[93][98] = 16'sd7;
        fc1_weights[93][99] = 16'sd67;
        fc1_weights[93][100] = 16'sd29;
        fc1_weights[93][101] = 16'sd-2;
        fc1_weights[93][102] = 16'sd58;
        fc1_weights[93][103] = 16'sd56;
        fc1_weights[93][104] = 16'sd-32;
        fc1_weights[93][105] = 16'sd-7;
        fc1_weights[93][106] = 16'sd2;
        fc1_weights[93][107] = 16'sd20;
        fc1_weights[93][108] = 16'sd8;
        fc1_weights[93][109] = 16'sd28;
        fc1_weights[93][110] = 16'sd4;
        fc1_weights[93][111] = 16'sd30;
        fc1_weights[93][112] = 16'sd0;
        fc1_weights[93][113] = 16'sd13;
        fc1_weights[93][114] = 16'sd20;
        fc1_weights[93][115] = 16'sd-24;
        fc1_weights[93][116] = 16'sd-31;
        fc1_weights[93][117] = 16'sd-27;
        fc1_weights[93][118] = 16'sd14;
        fc1_weights[93][119] = 16'sd80;
        fc1_weights[93][120] = 16'sd88;
        fc1_weights[93][121] = 16'sd-35;
        fc1_weights[93][122] = 16'sd-17;
        fc1_weights[93][123] = 16'sd27;
        fc1_weights[93][124] = 16'sd22;
        fc1_weights[93][125] = 16'sd100;
        fc1_weights[93][126] = 16'sd38;
        fc1_weights[93][127] = 16'sd14;
        fc1_weights[93][128] = 16'sd27;
        fc1_weights[93][129] = 16'sd123;
        fc1_weights[93][130] = 16'sd-44;
        fc1_weights[93][131] = 16'sd-58;
        fc1_weights[93][132] = 16'sd-42;
        fc1_weights[93][133] = 16'sd-58;
        fc1_weights[93][134] = 16'sd-1;
        fc1_weights[93][135] = 16'sd-39;
        fc1_weights[93][136] = 16'sd-48;
        fc1_weights[93][137] = 16'sd-12;
        fc1_weights[93][138] = 16'sd-121;
        fc1_weights[93][139] = 16'sd-58;
        fc1_weights[93][140] = 16'sd-4;
        fc1_weights[93][141] = 16'sd-17;
        fc1_weights[93][142] = 16'sd-67;
        fc1_weights[93][143] = 16'sd-37;
        fc1_weights[93][144] = 16'sd-36;
        fc1_weights[93][145] = 16'sd-18;
        fc1_weights[93][146] = 16'sd19;
        fc1_weights[93][147] = 16'sd-8;
        fc1_weights[93][148] = 16'sd41;
        fc1_weights[93][149] = 16'sd52;
        fc1_weights[93][150] = 16'sd43;
        fc1_weights[93][151] = 16'sd50;
        fc1_weights[93][152] = 16'sd25;
        fc1_weights[93][153] = 16'sd38;
        fc1_weights[93][154] = 16'sd32;
        fc1_weights[93][155] = 16'sd-15;
        fc1_weights[93][156] = 16'sd13;
        fc1_weights[93][157] = 16'sd4;
        fc1_weights[93][158] = 16'sd22;
        fc1_weights[93][159] = 16'sd3;
        fc1_weights[93][160] = 16'sd1;
        fc1_weights[93][161] = 16'sd51;
        fc1_weights[93][162] = 16'sd-25;
        fc1_weights[93][163] = 16'sd45;
        fc1_weights[93][164] = 16'sd-56;
        fc1_weights[93][165] = 16'sd13;
        fc1_weights[93][166] = 16'sd-90;
        fc1_weights[93][167] = 16'sd-68;
        fc1_weights[93][168] = 16'sd-93;
        fc1_weights[93][169] = 16'sd-41;
        fc1_weights[93][170] = 16'sd-46;
        fc1_weights[93][171] = 16'sd-44;
        fc1_weights[93][172] = 16'sd-29;
        fc1_weights[93][173] = 16'sd0;
        fc1_weights[93][174] = 16'sd16;
        fc1_weights[93][175] = 16'sd40;
        fc1_weights[93][176] = 16'sd51;
        fc1_weights[93][177] = 16'sd23;
        fc1_weights[93][178] = 16'sd63;
        fc1_weights[93][179] = 16'sd-3;
        fc1_weights[93][180] = 16'sd43;
        fc1_weights[93][181] = 16'sd-69;
        fc1_weights[93][182] = 16'sd-30;
        fc1_weights[93][183] = 16'sd-37;
        fc1_weights[93][184] = 16'sd-6;
        fc1_weights[93][185] = 16'sd-71;
        fc1_weights[93][186] = 16'sd-49;
        fc1_weights[93][187] = 16'sd7;
        fc1_weights[93][188] = 16'sd-11;
        fc1_weights[93][189] = 16'sd8;
        fc1_weights[93][190] = 16'sd-38;
        fc1_weights[93][191] = 16'sd-86;
        fc1_weights[93][192] = 16'sd-20;
        fc1_weights[93][193] = 16'sd-77;
        fc1_weights[93][194] = 16'sd-36;
        fc1_weights[93][195] = 16'sd-30;
        fc1_weights[93][196] = 16'sd23;
        fc1_weights[93][197] = 16'sd-71;
        fc1_weights[93][198] = 16'sd-23;
        fc1_weights[93][199] = 16'sd14;
        fc1_weights[93][200] = 16'sd-43;
        fc1_weights[93][201] = 16'sd21;
        fc1_weights[93][202] = 16'sd35;
        fc1_weights[93][203] = 16'sd17;
        fc1_weights[93][204] = 16'sd-34;
        fc1_weights[93][205] = 16'sd-28;
        fc1_weights[93][206] = 16'sd57;
        fc1_weights[93][207] = 16'sd-32;
        fc1_weights[94][0] = 16'sd30;
        fc1_weights[94][1] = 16'sd-46;
        fc1_weights[94][2] = 16'sd2;
        fc1_weights[94][3] = 16'sd-22;
        fc1_weights[94][4] = 16'sd23;
        fc1_weights[94][5] = 16'sd-45;
        fc1_weights[94][6] = 16'sd-11;
        fc1_weights[94][7] = 16'sd-37;
        fc1_weights[94][8] = 16'sd-29;
        fc1_weights[94][9] = 16'sd-12;
        fc1_weights[94][10] = 16'sd35;
        fc1_weights[94][11] = 16'sd23;
        fc1_weights[94][12] = 16'sd9;
        fc1_weights[94][13] = 16'sd8;
        fc1_weights[94][14] = 16'sd-33;
        fc1_weights[94][15] = 16'sd-19;
        fc1_weights[94][16] = 16'sd24;
        fc1_weights[94][17] = 16'sd-5;
        fc1_weights[94][18] = 16'sd-14;
        fc1_weights[94][19] = 16'sd85;
        fc1_weights[94][20] = 16'sd35;
        fc1_weights[94][21] = 16'sd19;
        fc1_weights[94][22] = 16'sd-8;
        fc1_weights[94][23] = 16'sd-9;
        fc1_weights[94][24] = 16'sd18;
        fc1_weights[94][25] = 16'sd25;
        fc1_weights[94][26] = 16'sd68;
        fc1_weights[94][27] = 16'sd36;
        fc1_weights[94][28] = 16'sd-40;
        fc1_weights[94][29] = 16'sd33;
        fc1_weights[94][30] = 16'sd-12;
        fc1_weights[94][31] = 16'sd-85;
        fc1_weights[94][32] = 16'sd-26;
        fc1_weights[94][33] = 16'sd41;
        fc1_weights[94][34] = 16'sd-37;
        fc1_weights[94][35] = 16'sd-17;
        fc1_weights[94][36] = 16'sd-54;
        fc1_weights[94][37] = 16'sd-43;
        fc1_weights[94][38] = 16'sd-34;
        fc1_weights[94][39] = 16'sd47;
        fc1_weights[94][40] = 16'sd-10;
        fc1_weights[94][41] = 16'sd28;
        fc1_weights[94][42] = 16'sd24;
        fc1_weights[94][43] = 16'sd123;
        fc1_weights[94][44] = 16'sd85;
        fc1_weights[94][45] = 16'sd74;
        fc1_weights[94][46] = 16'sd62;
        fc1_weights[94][47] = 16'sd45;
        fc1_weights[94][48] = 16'sd17;
        fc1_weights[94][49] = 16'sd-9;
        fc1_weights[94][50] = 16'sd4;
        fc1_weights[94][51] = 16'sd-9;
        fc1_weights[94][52] = 16'sd0;
        fc1_weights[94][53] = 16'sd21;
        fc1_weights[94][54] = 16'sd7;
        fc1_weights[94][55] = 16'sd0;
        fc1_weights[94][56] = 16'sd-24;
        fc1_weights[94][57] = 16'sd-22;
        fc1_weights[94][58] = 16'sd41;
        fc1_weights[94][59] = 16'sd-1;
        fc1_weights[94][60] = 16'sd-20;
        fc1_weights[94][61] = 16'sd45;
        fc1_weights[94][62] = 16'sd46;
        fc1_weights[94][63] = 16'sd6;
        fc1_weights[94][64] = 16'sd-35;
        fc1_weights[94][65] = 16'sd-15;
        fc1_weights[94][66] = 16'sd-49;
        fc1_weights[94][67] = 16'sd3;
        fc1_weights[94][68] = 16'sd96;
        fc1_weights[94][69] = 16'sd43;
        fc1_weights[94][70] = 16'sd-13;
        fc1_weights[94][71] = 16'sd12;
        fc1_weights[94][72] = 16'sd17;
        fc1_weights[94][73] = 16'sd-29;
        fc1_weights[94][74] = 16'sd-34;
        fc1_weights[94][75] = 16'sd-3;
        fc1_weights[94][76] = 16'sd-33;
        fc1_weights[94][77] = 16'sd-11;
        fc1_weights[94][78] = 16'sd73;
        fc1_weights[94][79] = 16'sd16;
        fc1_weights[94][80] = 16'sd31;
        fc1_weights[94][81] = 16'sd-9;
        fc1_weights[94][82] = 16'sd71;
        fc1_weights[94][83] = 16'sd-44;
        fc1_weights[94][84] = 16'sd7;
        fc1_weights[94][85] = 16'sd33;
        fc1_weights[94][86] = 16'sd2;
        fc1_weights[94][87] = 16'sd-31;
        fc1_weights[94][88] = 16'sd0;
        fc1_weights[94][89] = 16'sd-53;
        fc1_weights[94][90] = 16'sd-65;
        fc1_weights[94][91] = 16'sd-8;
        fc1_weights[94][92] = 16'sd-73;
        fc1_weights[94][93] = 16'sd-6;
        fc1_weights[94][94] = 16'sd64;
        fc1_weights[94][95] = 16'sd-10;
        fc1_weights[94][96] = 16'sd-44;
        fc1_weights[94][97] = 16'sd12;
        fc1_weights[94][98] = 16'sd-57;
        fc1_weights[94][99] = 16'sd-32;
        fc1_weights[94][100] = 16'sd-32;
        fc1_weights[94][101] = 16'sd-13;
        fc1_weights[94][102] = 16'sd15;
        fc1_weights[94][103] = 16'sd-19;
        fc1_weights[94][104] = 16'sd9;
        fc1_weights[94][105] = 16'sd86;
        fc1_weights[94][106] = 16'sd-33;
        fc1_weights[94][107] = 16'sd-25;
        fc1_weights[94][108] = 16'sd69;
        fc1_weights[94][109] = 16'sd-20;
        fc1_weights[94][110] = 16'sd49;
        fc1_weights[94][111] = 16'sd-27;
        fc1_weights[94][112] = 16'sd-36;
        fc1_weights[94][113] = 16'sd53;
        fc1_weights[94][114] = 16'sd11;
        fc1_weights[94][115] = 16'sd62;
        fc1_weights[94][116] = 16'sd3;
        fc1_weights[94][117] = 16'sd-21;
        fc1_weights[94][118] = 16'sd-28;
        fc1_weights[94][119] = 16'sd-64;
        fc1_weights[94][120] = 16'sd-32;
        fc1_weights[94][121] = 16'sd-31;
        fc1_weights[94][122] = 16'sd17;
        fc1_weights[94][123] = 16'sd-4;
        fc1_weights[94][124] = 16'sd-35;
        fc1_weights[94][125] = 16'sd-34;
        fc1_weights[94][126] = 16'sd-16;
        fc1_weights[94][127] = 16'sd1;
        fc1_weights[94][128] = 16'sd-42;
        fc1_weights[94][129] = 16'sd-38;
        fc1_weights[94][130] = 16'sd66;
        fc1_weights[94][131] = 16'sd-52;
        fc1_weights[94][132] = 16'sd-6;
        fc1_weights[94][133] = 16'sd-15;
        fc1_weights[94][134] = 16'sd7;
        fc1_weights[94][135] = 16'sd-56;
        fc1_weights[94][136] = 16'sd-18;
        fc1_weights[94][137] = 16'sd13;
        fc1_weights[94][138] = 16'sd86;
        fc1_weights[94][139] = 16'sd106;
        fc1_weights[94][140] = 16'sd71;
        fc1_weights[94][141] = 16'sd33;
        fc1_weights[94][142] = 16'sd-45;
        fc1_weights[94][143] = 16'sd-9;
        fc1_weights[94][144] = 16'sd-12;
        fc1_weights[94][145] = 16'sd-15;
        fc1_weights[94][146] = 16'sd-65;
        fc1_weights[94][147] = 16'sd-13;
        fc1_weights[94][148] = 16'sd5;
        fc1_weights[94][149] = 16'sd54;
        fc1_weights[94][150] = 16'sd-35;
        fc1_weights[94][151] = 16'sd3;
        fc1_weights[94][152] = 16'sd67;
        fc1_weights[94][153] = 16'sd12;
        fc1_weights[94][154] = 16'sd28;
        fc1_weights[94][155] = 16'sd37;
        fc1_weights[94][156] = 16'sd-21;
        fc1_weights[94][157] = 16'sd3;
        fc1_weights[94][158] = 16'sd54;
        fc1_weights[94][159] = 16'sd-5;
        fc1_weights[94][160] = 16'sd-4;
        fc1_weights[94][161] = 16'sd-5;
        fc1_weights[94][162] = 16'sd-68;
        fc1_weights[94][163] = 16'sd-20;
        fc1_weights[94][164] = 16'sd19;
        fc1_weights[94][165] = 16'sd36;
        fc1_weights[94][166] = 16'sd-14;
        fc1_weights[94][167] = 16'sd12;
        fc1_weights[94][168] = 16'sd-12;
        fc1_weights[94][169] = 16'sd6;
        fc1_weights[94][170] = 16'sd8;
        fc1_weights[94][171] = 16'sd30;
        fc1_weights[94][172] = 16'sd1;
        fc1_weights[94][173] = 16'sd35;
        fc1_weights[94][174] = 16'sd-40;
        fc1_weights[94][175] = 16'sd-16;
        fc1_weights[94][176] = 16'sd-13;
        fc1_weights[94][177] = 16'sd21;
        fc1_weights[94][178] = 16'sd22;
        fc1_weights[94][179] = 16'sd23;
        fc1_weights[94][180] = 16'sd-4;
        fc1_weights[94][181] = 16'sd-3;
        fc1_weights[94][182] = 16'sd37;
        fc1_weights[94][183] = 16'sd35;
        fc1_weights[94][184] = 16'sd36;
        fc1_weights[94][185] = 16'sd43;
        fc1_weights[94][186] = 16'sd-25;
        fc1_weights[94][187] = 16'sd18;
        fc1_weights[94][188] = 16'sd12;
        fc1_weights[94][189] = 16'sd-53;
        fc1_weights[94][190] = 16'sd-15;
        fc1_weights[94][191] = 16'sd-34;
        fc1_weights[94][192] = 16'sd-62;
        fc1_weights[94][193] = 16'sd-36;
        fc1_weights[94][194] = 16'sd-68;
        fc1_weights[94][195] = 16'sd-37;
        fc1_weights[94][196] = 16'sd-44;
        fc1_weights[94][197] = 16'sd-45;
        fc1_weights[94][198] = 16'sd29;
        fc1_weights[94][199] = 16'sd-58;
        fc1_weights[94][200] = 16'sd-32;
        fc1_weights[94][201] = 16'sd-30;
        fc1_weights[94][202] = 16'sd6;
        fc1_weights[94][203] = 16'sd-43;
        fc1_weights[94][204] = 16'sd13;
        fc1_weights[94][205] = 16'sd18;
        fc1_weights[94][206] = 16'sd-28;
        fc1_weights[94][207] = 16'sd-14;
        fc1_weights[95][0] = 16'sd22;
        fc1_weights[95][1] = 16'sd22;
        fc1_weights[95][2] = 16'sd-6;
        fc1_weights[95][3] = 16'sd13;
        fc1_weights[95][4] = 16'sd23;
        fc1_weights[95][5] = 16'sd5;
        fc1_weights[95][6] = 16'sd-3;
        fc1_weights[95][7] = 16'sd4;
        fc1_weights[95][8] = 16'sd32;
        fc1_weights[95][9] = 16'sd15;
        fc1_weights[95][10] = 16'sd8;
        fc1_weights[95][11] = 16'sd42;
        fc1_weights[95][12] = 16'sd-2;
        fc1_weights[95][13] = 16'sd5;
        fc1_weights[95][14] = 16'sd7;
        fc1_weights[95][15] = 16'sd15;
        fc1_weights[95][16] = 16'sd5;
        fc1_weights[95][17] = 16'sd-15;
        fc1_weights[95][18] = 16'sd-2;
        fc1_weights[95][19] = 16'sd-11;
        fc1_weights[95][20] = 16'sd-19;
        fc1_weights[95][21] = 16'sd-23;
        fc1_weights[95][22] = 16'sd-30;
        fc1_weights[95][23] = 16'sd20;
        fc1_weights[95][24] = 16'sd-2;
        fc1_weights[95][25] = 16'sd17;
        fc1_weights[95][26] = 16'sd-2;
        fc1_weights[95][27] = 16'sd20;
        fc1_weights[95][28] = 16'sd1;
        fc1_weights[95][29] = 16'sd15;
        fc1_weights[95][30] = 16'sd19;
        fc1_weights[95][31] = 16'sd3;
        fc1_weights[95][32] = 16'sd-2;
        fc1_weights[95][33] = 16'sd14;
        fc1_weights[95][34] = 16'sd9;
        fc1_weights[95][35] = 16'sd-13;
        fc1_weights[95][36] = 16'sd18;
        fc1_weights[95][37] = 16'sd25;
        fc1_weights[95][38] = 16'sd8;
        fc1_weights[95][39] = 16'sd51;
        fc1_weights[95][40] = 16'sd13;
        fc1_weights[95][41] = 16'sd8;
        fc1_weights[95][42] = 16'sd14;
        fc1_weights[95][43] = 16'sd18;
        fc1_weights[95][44] = 16'sd3;
        fc1_weights[95][45] = 16'sd-5;
        fc1_weights[95][46] = 16'sd-28;
        fc1_weights[95][47] = 16'sd-10;
        fc1_weights[95][48] = 16'sd-21;
        fc1_weights[95][49] = 16'sd-5;
        fc1_weights[95][50] = 16'sd-21;
        fc1_weights[95][51] = 16'sd-10;
        fc1_weights[95][52] = 16'sd2;
        fc1_weights[95][53] = 16'sd1;
        fc1_weights[95][54] = 16'sd-3;
        fc1_weights[95][55] = 16'sd-14;
        fc1_weights[95][56] = 16'sd3;
        fc1_weights[95][57] = 16'sd-19;
        fc1_weights[95][58] = 16'sd-31;
        fc1_weights[95][59] = 16'sd3;
        fc1_weights[95][60] = 16'sd-29;
        fc1_weights[95][61] = 16'sd-1;
        fc1_weights[95][62] = 16'sd3;
        fc1_weights[95][63] = 16'sd6;
        fc1_weights[95][64] = 16'sd7;
        fc1_weights[95][65] = 16'sd25;
        fc1_weights[95][66] = 16'sd20;
        fc1_weights[95][67] = 16'sd1;
        fc1_weights[95][68] = 16'sd-1;
        fc1_weights[95][69] = 16'sd2;
        fc1_weights[95][70] = 16'sd-11;
        fc1_weights[95][71] = 16'sd2;
        fc1_weights[95][72] = 16'sd-5;
        fc1_weights[95][73] = 16'sd1;
        fc1_weights[95][74] = 16'sd9;
        fc1_weights[95][75] = 16'sd9;
        fc1_weights[95][76] = 16'sd3;
        fc1_weights[95][77] = 16'sd-8;
        fc1_weights[95][78] = 16'sd22;
        fc1_weights[95][79] = 16'sd-17;
        fc1_weights[95][80] = 16'sd23;
        fc1_weights[95][81] = 16'sd12;
        fc1_weights[95][82] = 16'sd19;
        fc1_weights[95][83] = 16'sd33;
        fc1_weights[95][84] = 16'sd-27;
        fc1_weights[95][85] = 16'sd32;
        fc1_weights[95][86] = 16'sd9;
        fc1_weights[95][87] = 16'sd15;
        fc1_weights[95][88] = 16'sd24;
        fc1_weights[95][89] = 16'sd-5;
        fc1_weights[95][90] = 16'sd10;
        fc1_weights[95][91] = 16'sd-7;
        fc1_weights[95][92] = 16'sd-29;
        fc1_weights[95][93] = 16'sd-11;
        fc1_weights[95][94] = 16'sd-14;
        fc1_weights[95][95] = 16'sd0;
        fc1_weights[95][96] = 16'sd-7;
        fc1_weights[95][97] = 16'sd8;
        fc1_weights[95][98] = 16'sd-12;
        fc1_weights[95][99] = 16'sd-13;
        fc1_weights[95][100] = 16'sd1;
        fc1_weights[95][101] = 16'sd-7;
        fc1_weights[95][102] = 16'sd7;
        fc1_weights[95][103] = 16'sd2;
        fc1_weights[95][104] = 16'sd32;
        fc1_weights[95][105] = 16'sd29;
        fc1_weights[95][106] = 16'sd29;
        fc1_weights[95][107] = 16'sd23;
        fc1_weights[95][108] = 16'sd12;
        fc1_weights[95][109] = 16'sd30;
        fc1_weights[95][110] = 16'sd26;
        fc1_weights[95][111] = 16'sd88;
        fc1_weights[95][112] = 16'sd75;
        fc1_weights[95][113] = 16'sd38;
        fc1_weights[95][114] = 16'sd38;
        fc1_weights[95][115] = 16'sd-3;
        fc1_weights[95][116] = 16'sd-13;
        fc1_weights[95][117] = 16'sd-37;
        fc1_weights[95][118] = 16'sd-5;
        fc1_weights[95][119] = 16'sd-42;
        fc1_weights[95][120] = 16'sd-26;
        fc1_weights[95][121] = 16'sd-9;
        fc1_weights[95][122] = 16'sd8;
        fc1_weights[95][123] = 16'sd26;
        fc1_weights[95][124] = 16'sd3;
        fc1_weights[95][125] = 16'sd-8;
        fc1_weights[95][126] = 16'sd7;
        fc1_weights[95][127] = 16'sd19;
        fc1_weights[95][128] = 16'sd21;
        fc1_weights[95][129] = 16'sd-4;
        fc1_weights[95][130] = 16'sd33;
        fc1_weights[95][131] = 16'sd26;
        fc1_weights[95][132] = 16'sd21;
        fc1_weights[95][133] = 16'sd13;
        fc1_weights[95][134] = 16'sd34;
        fc1_weights[95][135] = 16'sd41;
        fc1_weights[95][136] = 16'sd17;
        fc1_weights[95][137] = 16'sd36;
        fc1_weights[95][138] = 16'sd22;
        fc1_weights[95][139] = 16'sd17;
        fc1_weights[95][140] = 16'sd23;
        fc1_weights[95][141] = 16'sd26;
        fc1_weights[95][142] = 16'sd25;
        fc1_weights[95][143] = 16'sd22;
        fc1_weights[95][144] = 16'sd12;
        fc1_weights[95][145] = 16'sd-1;
        fc1_weights[95][146] = 16'sd-15;
        fc1_weights[95][147] = 16'sd-16;
        fc1_weights[95][148] = 16'sd7;
        fc1_weights[95][149] = 16'sd-22;
        fc1_weights[95][150] = 16'sd7;
        fc1_weights[95][151] = 16'sd-21;
        fc1_weights[95][152] = 16'sd-25;
        fc1_weights[95][153] = 16'sd-18;
        fc1_weights[95][154] = 16'sd-20;
        fc1_weights[95][155] = 16'sd-10;
        fc1_weights[95][156] = 16'sd33;
        fc1_weights[95][157] = 16'sd22;
        fc1_weights[95][158] = 16'sd-6;
        fc1_weights[95][159] = 16'sd6;
        fc1_weights[95][160] = 16'sd6;
        fc1_weights[95][161] = 16'sd-14;
        fc1_weights[95][162] = 16'sd29;
        fc1_weights[95][163] = 16'sd14;
        fc1_weights[95][164] = 16'sd17;
        fc1_weights[95][165] = 16'sd-10;
        fc1_weights[95][166] = 16'sd-15;
        fc1_weights[95][167] = 16'sd-16;
        fc1_weights[95][168] = 16'sd7;
        fc1_weights[95][169] = 16'sd25;
        fc1_weights[95][170] = 16'sd25;
        fc1_weights[95][171] = 16'sd36;
        fc1_weights[95][172] = 16'sd11;
        fc1_weights[95][173] = 16'sd-25;
        fc1_weights[95][174] = 16'sd-10;
        fc1_weights[95][175] = 16'sd-2;
        fc1_weights[95][176] = 16'sd-31;
        fc1_weights[95][177] = 16'sd-27;
        fc1_weights[95][178] = 16'sd-37;
        fc1_weights[95][179] = 16'sd-17;
        fc1_weights[95][180] = 16'sd-12;
        fc1_weights[95][181] = 16'sd-22;
        fc1_weights[95][182] = 16'sd2;
        fc1_weights[95][183] = 16'sd-8;
        fc1_weights[95][184] = 16'sd-18;
        fc1_weights[95][185] = 16'sd-6;
        fc1_weights[95][186] = 16'sd24;
        fc1_weights[95][187] = 16'sd9;
        fc1_weights[95][188] = 16'sd16;
        fc1_weights[95][189] = 16'sd29;
        fc1_weights[95][190] = 16'sd-6;
        fc1_weights[95][191] = 16'sd-11;
        fc1_weights[95][192] = 16'sd0;
        fc1_weights[95][193] = 16'sd2;
        fc1_weights[95][194] = 16'sd8;
        fc1_weights[95][195] = 16'sd-11;
        fc1_weights[95][196] = 16'sd8;
        fc1_weights[95][197] = 16'sd12;
        fc1_weights[95][198] = 16'sd33;
        fc1_weights[95][199] = 16'sd4;
        fc1_weights[95][200] = 16'sd-2;
        fc1_weights[95][201] = 16'sd0;
        fc1_weights[95][202] = 16'sd-11;
        fc1_weights[95][203] = 16'sd10;
        fc1_weights[95][204] = 16'sd14;
        fc1_weights[95][205] = 16'sd-37;
        fc1_weights[95][206] = 16'sd-16;
        fc1_weights[95][207] = 16'sd-22;
        fc1_weights[96][0] = 16'sd-25;
        fc1_weights[96][1] = 16'sd-13;
        fc1_weights[96][2] = 16'sd-36;
        fc1_weights[96][3] = 16'sd-15;
        fc1_weights[96][4] = 16'sd-44;
        fc1_weights[96][5] = 16'sd6;
        fc1_weights[96][6] = 16'sd26;
        fc1_weights[96][7] = 16'sd-7;
        fc1_weights[96][8] = 16'sd4;
        fc1_weights[96][9] = 16'sd29;
        fc1_weights[96][10] = 16'sd36;
        fc1_weights[96][11] = 16'sd-51;
        fc1_weights[96][12] = 16'sd-87;
        fc1_weights[96][13] = 16'sd-97;
        fc1_weights[96][14] = 16'sd-58;
        fc1_weights[96][15] = 16'sd30;
        fc1_weights[96][16] = 16'sd45;
        fc1_weights[96][17] = 16'sd-11;
        fc1_weights[96][18] = 16'sd-30;
        fc1_weights[96][19] = 16'sd-29;
        fc1_weights[96][20] = 16'sd15;
        fc1_weights[96][21] = 16'sd-49;
        fc1_weights[96][22] = 16'sd-29;
        fc1_weights[96][23] = 16'sd-44;
        fc1_weights[96][24] = 16'sd54;
        fc1_weights[96][25] = 16'sd7;
        fc1_weights[96][26] = 16'sd-64;
        fc1_weights[96][27] = 16'sd-70;
        fc1_weights[96][28] = 16'sd-56;
        fc1_weights[96][29] = 16'sd-41;
        fc1_weights[96][30] = 16'sd27;
        fc1_weights[96][31] = 16'sd26;
        fc1_weights[96][32] = 16'sd12;
        fc1_weights[96][33] = 16'sd-45;
        fc1_weights[96][34] = 16'sd33;
        fc1_weights[96][35] = 16'sd5;
        fc1_weights[96][36] = 16'sd18;
        fc1_weights[96][37] = 16'sd48;
        fc1_weights[96][38] = 16'sd-36;
        fc1_weights[96][39] = 16'sd-127;
        fc1_weights[96][40] = 16'sd96;
        fc1_weights[96][41] = 16'sd81;
        fc1_weights[96][42] = 16'sd-15;
        fc1_weights[96][43] = 16'sd-21;
        fc1_weights[96][44] = 16'sd-18;
        fc1_weights[96][45] = 16'sd-99;
        fc1_weights[96][46] = 16'sd-6;
        fc1_weights[96][47] = 16'sd-65;
        fc1_weights[96][48] = 16'sd25;
        fc1_weights[96][49] = 16'sd34;
        fc1_weights[96][50] = 16'sd-13;
        fc1_weights[96][51] = 16'sd-35;
        fc1_weights[96][52] = 16'sd-107;
        fc1_weights[96][53] = 16'sd-35;
        fc1_weights[96][54] = 16'sd47;
        fc1_weights[96][55] = 16'sd5;
        fc1_weights[96][56] = 16'sd12;
        fc1_weights[96][57] = 16'sd10;
        fc1_weights[96][58] = 16'sd-15;
        fc1_weights[96][59] = 16'sd-50;
        fc1_weights[96][60] = 16'sd18;
        fc1_weights[96][61] = 16'sd-34;
        fc1_weights[96][62] = 16'sd-54;
        fc1_weights[96][63] = 16'sd0;
        fc1_weights[96][64] = 16'sd-16;
        fc1_weights[96][65] = 16'sd3;
        fc1_weights[96][66] = 16'sd33;
        fc1_weights[96][67] = 16'sd-12;
        fc1_weights[96][68] = 16'sd-22;
        fc1_weights[96][69] = 16'sd-28;
        fc1_weights[96][70] = 16'sd-69;
        fc1_weights[96][71] = 16'sd-10;
        fc1_weights[96][72] = 16'sd2;
        fc1_weights[96][73] = 16'sd-59;
        fc1_weights[96][74] = 16'sd-15;
        fc1_weights[96][75] = 16'sd-7;
        fc1_weights[96][76] = 16'sd7;
        fc1_weights[96][77] = 16'sd-28;
        fc1_weights[96][78] = 16'sd-2;
        fc1_weights[96][79] = 16'sd71;
        fc1_weights[96][80] = 16'sd1;
        fc1_weights[96][81] = 16'sd8;
        fc1_weights[96][82] = 16'sd26;
        fc1_weights[96][83] = 16'sd20;
        fc1_weights[96][84] = 16'sd0;
        fc1_weights[96][85] = 16'sd-43;
        fc1_weights[96][86] = 16'sd19;
        fc1_weights[96][87] = 16'sd-37;
        fc1_weights[96][88] = 16'sd-59;
        fc1_weights[96][89] = 16'sd103;
        fc1_weights[96][90] = 16'sd8;
        fc1_weights[96][91] = 16'sd32;
        fc1_weights[96][92] = 16'sd38;
        fc1_weights[96][93] = 16'sd91;
        fc1_weights[96][94] = 16'sd24;
        fc1_weights[96][95] = 16'sd18;
        fc1_weights[96][96] = 16'sd-2;
        fc1_weights[96][97] = 16'sd7;
        fc1_weights[96][98] = 16'sd-1;
        fc1_weights[96][99] = 16'sd-5;
        fc1_weights[96][100] = 16'sd30;
        fc1_weights[96][101] = 16'sd-13;
        fc1_weights[96][102] = 16'sd-4;
        fc1_weights[96][103] = 16'sd-79;
        fc1_weights[96][104] = 16'sd7;
        fc1_weights[96][105] = 16'sd-24;
        fc1_weights[96][106] = 16'sd-13;
        fc1_weights[96][107] = 16'sd-32;
        fc1_weights[96][108] = 16'sd34;
        fc1_weights[96][109] = 16'sd-24;
        fc1_weights[96][110] = 16'sd24;
        fc1_weights[96][111] = 16'sd-48;
        fc1_weights[96][112] = 16'sd69;
        fc1_weights[96][113] = 16'sd58;
        fc1_weights[96][114] = 16'sd19;
        fc1_weights[96][115] = 16'sd-27;
        fc1_weights[96][116] = 16'sd29;
        fc1_weights[96][117] = 16'sd45;
        fc1_weights[96][118] = 16'sd25;
        fc1_weights[96][119] = 16'sd30;
        fc1_weights[96][120] = 16'sd29;
        fc1_weights[96][121] = 16'sd61;
        fc1_weights[96][122] = 16'sd90;
        fc1_weights[96][123] = 16'sd22;
        fc1_weights[96][124] = 16'sd-65;
        fc1_weights[96][125] = 16'sd-19;
        fc1_weights[96][126] = 16'sd-58;
        fc1_weights[96][127] = 16'sd-37;
        fc1_weights[96][128] = 16'sd-40;
        fc1_weights[96][129] = 16'sd-105;
        fc1_weights[96][130] = 16'sd-19;
        fc1_weights[96][131] = 16'sd-53;
        fc1_weights[96][132] = 16'sd49;
        fc1_weights[96][133] = 16'sd11;
        fc1_weights[96][134] = 16'sd58;
        fc1_weights[96][135] = 16'sd48;
        fc1_weights[96][136] = 16'sd-54;
        fc1_weights[96][137] = 16'sd1;
        fc1_weights[96][138] = 16'sd-8;
        fc1_weights[96][139] = 16'sd61;
        fc1_weights[96][140] = 16'sd85;
        fc1_weights[96][141] = 16'sd-57;
        fc1_weights[96][142] = 16'sd45;
        fc1_weights[96][143] = 16'sd19;
        fc1_weights[96][144] = 16'sd70;
        fc1_weights[96][145] = 16'sd-10;
        fc1_weights[96][146] = 16'sd-7;
        fc1_weights[96][147] = 16'sd11;
        fc1_weights[96][148] = 16'sd33;
        fc1_weights[96][149] = 16'sd-21;
        fc1_weights[96][150] = 16'sd-19;
        fc1_weights[96][151] = 16'sd-43;
        fc1_weights[96][152] = 16'sd-53;
        fc1_weights[96][153] = 16'sd-24;
        fc1_weights[96][154] = 16'sd-31;
        fc1_weights[96][155] = 16'sd34;
        fc1_weights[96][156] = 16'sd33;
        fc1_weights[96][157] = 16'sd29;
        fc1_weights[96][158] = 16'sd-10;
        fc1_weights[96][159] = 16'sd15;
        fc1_weights[96][160] = 16'sd-58;
        fc1_weights[96][161] = 16'sd-111;
        fc1_weights[96][162] = 16'sd-44;
        fc1_weights[96][163] = 16'sd-1;
        fc1_weights[96][164] = 16'sd51;
        fc1_weights[96][165] = 16'sd74;
        fc1_weights[96][166] = 16'sd74;
        fc1_weights[96][167] = 16'sd27;
        fc1_weights[96][168] = 16'sd75;
        fc1_weights[96][169] = 16'sd-15;
        fc1_weights[96][170] = 16'sd-27;
        fc1_weights[96][171] = 16'sd44;
        fc1_weights[96][172] = 16'sd44;
        fc1_weights[96][173] = 16'sd59;
        fc1_weights[96][174] = 16'sd-29;
        fc1_weights[96][175] = 16'sd10;
        fc1_weights[96][176] = 16'sd0;
        fc1_weights[96][177] = 16'sd32;
        fc1_weights[96][178] = 16'sd-52;
        fc1_weights[96][179] = 16'sd-4;
        fc1_weights[96][180] = 16'sd38;
        fc1_weights[96][181] = 16'sd3;
        fc1_weights[96][182] = 16'sd-10;
        fc1_weights[96][183] = 16'sd-14;
        fc1_weights[96][184] = 16'sd-41;
        fc1_weights[96][185] = 16'sd94;
        fc1_weights[96][186] = 16'sd-42;
        fc1_weights[96][187] = 16'sd40;
        fc1_weights[96][188] = 16'sd18;
        fc1_weights[96][189] = 16'sd-5;
        fc1_weights[96][190] = 16'sd54;
        fc1_weights[96][191] = 16'sd99;
        fc1_weights[96][192] = 16'sd-13;
        fc1_weights[96][193] = 16'sd17;
        fc1_weights[96][194] = 16'sd9;
        fc1_weights[96][195] = 16'sd-20;
        fc1_weights[96][196] = 16'sd-28;
        fc1_weights[96][197] = 16'sd50;
        fc1_weights[96][198] = 16'sd15;
        fc1_weights[96][199] = 16'sd71;
        fc1_weights[96][200] = 16'sd-40;
        fc1_weights[96][201] = 16'sd-4;
        fc1_weights[96][202] = 16'sd-17;
        fc1_weights[96][203] = 16'sd70;
        fc1_weights[96][204] = 16'sd-13;
        fc1_weights[96][205] = 16'sd46;
        fc1_weights[96][206] = 16'sd3;
        fc1_weights[96][207] = 16'sd-52;
        fc1_weights[97][0] = 16'sd-6;
        fc1_weights[97][1] = 16'sd-12;
        fc1_weights[97][2] = 16'sd6;
        fc1_weights[97][3] = 16'sd-10;
        fc1_weights[97][4] = 16'sd-49;
        fc1_weights[97][5] = 16'sd14;
        fc1_weights[97][6] = 16'sd-88;
        fc1_weights[97][7] = 16'sd-7;
        fc1_weights[97][8] = 16'sd-45;
        fc1_weights[97][9] = 16'sd-9;
        fc1_weights[97][10] = 16'sd69;
        fc1_weights[97][11] = 16'sd43;
        fc1_weights[97][12] = 16'sd70;
        fc1_weights[97][13] = 16'sd111;
        fc1_weights[97][14] = 16'sd42;
        fc1_weights[97][15] = 16'sd-14;
        fc1_weights[97][16] = 16'sd-4;
        fc1_weights[97][17] = 16'sd-26;
        fc1_weights[97][18] = 16'sd-9;
        fc1_weights[97][19] = 16'sd6;
        fc1_weights[97][20] = 16'sd-37;
        fc1_weights[97][21] = 16'sd57;
        fc1_weights[97][22] = 16'sd42;
        fc1_weights[97][23] = 16'sd104;
        fc1_weights[97][24] = 16'sd38;
        fc1_weights[97][25] = 16'sd48;
        fc1_weights[97][26] = 16'sd-16;
        fc1_weights[97][27] = 16'sd-51;
        fc1_weights[97][28] = 16'sd27;
        fc1_weights[97][29] = 16'sd49;
        fc1_weights[97][30] = 16'sd-1;
        fc1_weights[97][31] = 16'sd2;
        fc1_weights[97][32] = 16'sd-44;
        fc1_weights[97][33] = 16'sd-82;
        fc1_weights[97][34] = 16'sd-31;
        fc1_weights[97][35] = 16'sd-68;
        fc1_weights[97][36] = 16'sd39;
        fc1_weights[97][37] = 16'sd103;
        fc1_weights[97][38] = 16'sd61;
        fc1_weights[97][39] = 16'sd57;
        fc1_weights[97][40] = 16'sd-3;
        fc1_weights[97][41] = 16'sd-55;
        fc1_weights[97][42] = 16'sd11;
        fc1_weights[97][43] = 16'sd-88;
        fc1_weights[97][44] = 16'sd-16;
        fc1_weights[97][45] = 16'sd-16;
        fc1_weights[97][46] = 16'sd-9;
        fc1_weights[97][47] = 16'sd2;
        fc1_weights[97][48] = 16'sd-17;
        fc1_weights[97][49] = 16'sd-33;
        fc1_weights[97][50] = 16'sd32;
        fc1_weights[97][51] = 16'sd-30;
        fc1_weights[97][52] = 16'sd52;
        fc1_weights[97][53] = 16'sd15;
        fc1_weights[97][54] = 16'sd-3;
        fc1_weights[97][55] = 16'sd52;
        fc1_weights[97][56] = 16'sd39;
        fc1_weights[97][57] = 16'sd24;
        fc1_weights[97][58] = 16'sd-10;
        fc1_weights[97][59] = 16'sd-9;
        fc1_weights[97][60] = 16'sd-42;
        fc1_weights[97][61] = 16'sd-73;
        fc1_weights[97][62] = 16'sd-86;
        fc1_weights[97][63] = 16'sd-6;
        fc1_weights[97][64] = 16'sd47;
        fc1_weights[97][65] = 16'sd-3;
        fc1_weights[97][66] = 16'sd14;
        fc1_weights[97][67] = 16'sd-19;
        fc1_weights[97][68] = 16'sd-63;
        fc1_weights[97][69] = 16'sd-2;
        fc1_weights[97][70] = 16'sd21;
        fc1_weights[97][71] = 16'sd-72;
        fc1_weights[97][72] = 16'sd-86;
        fc1_weights[97][73] = 16'sd-2;
        fc1_weights[97][74] = 16'sd-10;
        fc1_weights[97][75] = 16'sd3;
        fc1_weights[97][76] = 16'sd10;
        fc1_weights[97][77] = 16'sd29;
        fc1_weights[97][78] = 16'sd-30;
        fc1_weights[97][79] = 16'sd-88;
        fc1_weights[97][80] = 16'sd9;
        fc1_weights[97][81] = 16'sd11;
        fc1_weights[97][82] = 16'sd18;
        fc1_weights[97][83] = 16'sd74;
        fc1_weights[97][84] = 16'sd9;
        fc1_weights[97][85] = 16'sd33;
        fc1_weights[97][86] = 16'sd18;
        fc1_weights[97][87] = 16'sd41;
        fc1_weights[97][88] = 16'sd-35;
        fc1_weights[97][89] = 16'sd-64;
        fc1_weights[97][90] = 16'sd13;
        fc1_weights[97][91] = 16'sd-39;
        fc1_weights[97][92] = 16'sd-36;
        fc1_weights[97][93] = 16'sd-33;
        fc1_weights[97][94] = 16'sd-43;
        fc1_weights[97][95] = 16'sd33;
        fc1_weights[97][96] = 16'sd-22;
        fc1_weights[97][97] = 16'sd10;
        fc1_weights[97][98] = 16'sd-4;
        fc1_weights[97][99] = 16'sd12;
        fc1_weights[97][100] = 16'sd-31;
        fc1_weights[97][101] = 16'sd-4;
        fc1_weights[97][102] = 16'sd-28;
        fc1_weights[97][103] = 16'sd7;
        fc1_weights[97][104] = 16'sd-7;
        fc1_weights[97][105] = 16'sd-24;
        fc1_weights[97][106] = 16'sd44;
        fc1_weights[97][107] = 16'sd0;
        fc1_weights[97][108] = 16'sd-16;
        fc1_weights[97][109] = 16'sd35;
        fc1_weights[97][110] = 16'sd-39;
        fc1_weights[97][111] = 16'sd76;
        fc1_weights[97][112] = 16'sd59;
        fc1_weights[97][113] = 16'sd-42;
        fc1_weights[97][114] = 16'sd38;
        fc1_weights[97][115] = 16'sd29;
        fc1_weights[97][116] = 16'sd-53;
        fc1_weights[97][117] = 16'sd-37;
        fc1_weights[97][118] = 16'sd4;
        fc1_weights[97][119] = 16'sd-43;
        fc1_weights[97][120] = 16'sd37;
        fc1_weights[97][121] = 16'sd34;
        fc1_weights[97][122] = 16'sd25;
        fc1_weights[97][123] = 16'sd-30;
        fc1_weights[97][124] = 16'sd9;
        fc1_weights[97][125] = 16'sd-29;
        fc1_weights[97][126] = 16'sd42;
        fc1_weights[97][127] = 16'sd58;
        fc1_weights[97][128] = 16'sd-15;
        fc1_weights[97][129] = 16'sd77;
        fc1_weights[97][130] = 16'sd-66;
        fc1_weights[97][131] = 16'sd-49;
        fc1_weights[97][132] = 16'sd-24;
        fc1_weights[97][133] = 16'sd-37;
        fc1_weights[97][134] = 16'sd-37;
        fc1_weights[97][135] = 16'sd-9;
        fc1_weights[97][136] = 16'sd6;
        fc1_weights[97][137] = 16'sd-28;
        fc1_weights[97][138] = 16'sd56;
        fc1_weights[97][139] = 16'sd-14;
        fc1_weights[97][140] = 16'sd-34;
        fc1_weights[97][141] = 16'sd71;
        fc1_weights[97][142] = 16'sd13;
        fc1_weights[97][143] = 16'sd58;
        fc1_weights[97][144] = 16'sd-8;
        fc1_weights[97][145] = 16'sd38;
        fc1_weights[97][146] = 16'sd56;
        fc1_weights[97][147] = 16'sd3;
        fc1_weights[97][148] = 16'sd3;
        fc1_weights[97][149] = 16'sd-34;
        fc1_weights[97][150] = 16'sd52;
        fc1_weights[97][151] = 16'sd27;
        fc1_weights[97][152] = 16'sd19;
        fc1_weights[97][153] = 16'sd-53;
        fc1_weights[97][154] = 16'sd21;
        fc1_weights[97][155] = 16'sd38;
        fc1_weights[97][156] = 16'sd-74;
        fc1_weights[97][157] = 16'sd-45;
        fc1_weights[97][158] = 16'sd-57;
        fc1_weights[97][159] = 16'sd-84;
        fc1_weights[97][160] = 16'sd25;
        fc1_weights[97][161] = 16'sd83;
        fc1_weights[97][162] = 16'sd79;
        fc1_weights[97][163] = 16'sd25;
        fc1_weights[97][164] = 16'sd-1;
        fc1_weights[97][165] = 16'sd16;
        fc1_weights[97][166] = 16'sd-5;
        fc1_weights[97][167] = 16'sd-36;
        fc1_weights[97][168] = 16'sd-53;
        fc1_weights[97][169] = 16'sd-30;
        fc1_weights[97][170] = 16'sd-10;
        fc1_weights[97][171] = 16'sd-38;
        fc1_weights[97][172] = 16'sd30;
        fc1_weights[97][173] = 16'sd0;
        fc1_weights[97][174] = 16'sd7;
        fc1_weights[97][175] = 16'sd-25;
        fc1_weights[97][176] = 16'sd22;
        fc1_weights[97][177] = 16'sd18;
        fc1_weights[97][178] = 16'sd18;
        fc1_weights[97][179] = 16'sd46;
        fc1_weights[97][180] = 16'sd7;
        fc1_weights[97][181] = 16'sd38;
        fc1_weights[97][182] = 16'sd29;
        fc1_weights[97][183] = 16'sd-78;
        fc1_weights[97][184] = 16'sd-21;
        fc1_weights[97][185] = 16'sd-78;
        fc1_weights[97][186] = 16'sd62;
        fc1_weights[97][187] = 16'sd-9;
        fc1_weights[97][188] = 16'sd-1;
        fc1_weights[97][189] = 16'sd29;
        fc1_weights[97][190] = 16'sd-20;
        fc1_weights[97][191] = 16'sd-43;
        fc1_weights[97][192] = 16'sd38;
        fc1_weights[97][193] = 16'sd7;
        fc1_weights[97][194] = 16'sd-7;
        fc1_weights[97][195] = 16'sd35;
        fc1_weights[97][196] = 16'sd23;
        fc1_weights[97][197] = 16'sd26;
        fc1_weights[97][198] = 16'sd-34;
        fc1_weights[97][199] = 16'sd16;
        fc1_weights[97][200] = 16'sd48;
        fc1_weights[97][201] = 16'sd-42;
        fc1_weights[97][202] = 16'sd-43;
        fc1_weights[97][203] = 16'sd53;
        fc1_weights[97][204] = 16'sd34;
        fc1_weights[97][205] = 16'sd-16;
        fc1_weights[97][206] = 16'sd19;
        fc1_weights[97][207] = 16'sd60;
        fc1_weights[98][0] = 16'sd-3;
        fc1_weights[98][1] = 16'sd34;
        fc1_weights[98][2] = 16'sd-3;
        fc1_weights[98][3] = 16'sd-76;
        fc1_weights[98][4] = 16'sd-44;
        fc1_weights[98][5] = 16'sd-3;
        fc1_weights[98][6] = 16'sd31;
        fc1_weights[98][7] = 16'sd20;
        fc1_weights[98][8] = 16'sd-20;
        fc1_weights[98][9] = 16'sd-21;
        fc1_weights[98][10] = 16'sd-5;
        fc1_weights[98][11] = 16'sd-125;
        fc1_weights[98][12] = 16'sd-125;
        fc1_weights[98][13] = 16'sd-12;
        fc1_weights[98][14] = 16'sd-1;
        fc1_weights[98][15] = 16'sd25;
        fc1_weights[98][16] = 16'sd22;
        fc1_weights[98][17] = 16'sd6;
        fc1_weights[98][18] = 16'sd37;
        fc1_weights[98][19] = 16'sd-2;
        fc1_weights[98][20] = 16'sd36;
        fc1_weights[98][21] = 16'sd6;
        fc1_weights[98][22] = 16'sd37;
        fc1_weights[98][23] = 16'sd41;
        fc1_weights[98][24] = 16'sd36;
        fc1_weights[98][25] = 16'sd76;
        fc1_weights[98][26] = 16'sd24;
        fc1_weights[98][27] = 16'sd12;
        fc1_weights[98][28] = 16'sd30;
        fc1_weights[98][29] = 16'sd-2;
        fc1_weights[98][30] = 16'sd-49;
        fc1_weights[98][31] = 16'sd1;
        fc1_weights[98][32] = 16'sd-21;
        fc1_weights[98][33] = 16'sd-58;
        fc1_weights[98][34] = 16'sd-28;
        fc1_weights[98][35] = 16'sd39;
        fc1_weights[98][36] = 16'sd10;
        fc1_weights[98][37] = 16'sd-59;
        fc1_weights[98][38] = 16'sd-20;
        fc1_weights[98][39] = 16'sd-108;
        fc1_weights[98][40] = 16'sd27;
        fc1_weights[98][41] = 16'sd52;
        fc1_weights[98][42] = 16'sd-34;
        fc1_weights[98][43] = 16'sd-13;
        fc1_weights[98][44] = 16'sd13;
        fc1_weights[98][45] = 16'sd-41;
        fc1_weights[98][46] = 16'sd-6;
        fc1_weights[98][47] = 16'sd-36;
        fc1_weights[98][48] = 16'sd-13;
        fc1_weights[98][49] = 16'sd42;
        fc1_weights[98][50] = 16'sd34;
        fc1_weights[98][51] = 16'sd-23;
        fc1_weights[98][52] = 16'sd37;
        fc1_weights[98][53] = 16'sd22;
        fc1_weights[98][54] = 16'sd15;
        fc1_weights[98][55] = 16'sd15;
        fc1_weights[98][56] = 16'sd41;
        fc1_weights[98][57] = 16'sd42;
        fc1_weights[98][58] = 16'sd-7;
        fc1_weights[98][59] = 16'sd-48;
        fc1_weights[98][60] = 16'sd-7;
        fc1_weights[98][61] = 16'sd-23;
        fc1_weights[98][62] = 16'sd9;
        fc1_weights[98][63] = 16'sd42;
        fc1_weights[98][64] = 16'sd-9;
        fc1_weights[98][65] = 16'sd-42;
        fc1_weights[98][66] = 16'sd-18;
        fc1_weights[98][67] = 16'sd23;
        fc1_weights[98][68] = 16'sd-24;
        fc1_weights[98][69] = 16'sd29;
        fc1_weights[98][70] = 16'sd73;
        fc1_weights[98][71] = 16'sd6;
        fc1_weights[98][72] = 16'sd-46;
        fc1_weights[98][73] = 16'sd-50;
        fc1_weights[98][74] = 16'sd-39;
        fc1_weights[98][75] = 16'sd19;
        fc1_weights[98][76] = 16'sd24;
        fc1_weights[98][77] = 16'sd-13;
        fc1_weights[98][78] = 16'sd12;
        fc1_weights[98][79] = 16'sd35;
        fc1_weights[98][80] = 16'sd20;
        fc1_weights[98][81] = 16'sd26;
        fc1_weights[98][82] = 16'sd-48;
        fc1_weights[98][83] = 16'sd20;
        fc1_weights[98][84] = 16'sd-43;
        fc1_weights[98][85] = 16'sd-9;
        fc1_weights[98][86] = 16'sd-12;
        fc1_weights[98][87] = 16'sd-57;
        fc1_weights[98][88] = 16'sd-8;
        fc1_weights[98][89] = 16'sd27;
        fc1_weights[98][90] = 16'sd-85;
        fc1_weights[98][91] = 16'sd12;
        fc1_weights[98][92] = 16'sd-24;
        fc1_weights[98][93] = 16'sd-1;
        fc1_weights[98][94] = 16'sd-20;
        fc1_weights[98][95] = 16'sd-27;
        fc1_weights[98][96] = 16'sd42;
        fc1_weights[98][97] = 16'sd33;
        fc1_weights[98][98] = 16'sd40;
        fc1_weights[98][99] = 16'sd-20;
        fc1_weights[98][100] = 16'sd-23;
        fc1_weights[98][101] = 16'sd17;
        fc1_weights[98][102] = 16'sd19;
        fc1_weights[98][103] = 16'sd-52;
        fc1_weights[98][104] = 16'sd31;
        fc1_weights[98][105] = 16'sd10;
        fc1_weights[98][106] = 16'sd18;
        fc1_weights[98][107] = 16'sd-10;
        fc1_weights[98][108] = 16'sd-1;
        fc1_weights[98][109] = 16'sd48;
        fc1_weights[98][110] = 16'sd-53;
        fc1_weights[98][111] = 16'sd-23;
        fc1_weights[98][112] = 16'sd49;
        fc1_weights[98][113] = 16'sd-58;
        fc1_weights[98][114] = 16'sd9;
        fc1_weights[98][115] = 16'sd-13;
        fc1_weights[98][116] = 16'sd-37;
        fc1_weights[98][117] = 16'sd-9;
        fc1_weights[98][118] = 16'sd26;
        fc1_weights[98][119] = 16'sd-26;
        fc1_weights[98][120] = 16'sd-39;
        fc1_weights[98][121] = 16'sd-25;
        fc1_weights[98][122] = 16'sd-2;
        fc1_weights[98][123] = 16'sd16;
        fc1_weights[98][124] = 16'sd-52;
        fc1_weights[98][125] = 16'sd-55;
        fc1_weights[98][126] = 16'sd-57;
        fc1_weights[98][127] = 16'sd26;
        fc1_weights[98][128] = 16'sd-4;
        fc1_weights[98][129] = 16'sd6;
        fc1_weights[98][130] = 16'sd-53;
        fc1_weights[98][131] = 16'sd24;
        fc1_weights[98][132] = 16'sd8;
        fc1_weights[98][133] = 16'sd23;
        fc1_weights[98][134] = 16'sd6;
        fc1_weights[98][135] = 16'sd37;
        fc1_weights[98][136] = 16'sd22;
        fc1_weights[98][137] = 16'sd2;
        fc1_weights[98][138] = 16'sd28;
        fc1_weights[98][139] = 16'sd-75;
        fc1_weights[98][140] = 16'sd-53;
        fc1_weights[98][141] = 16'sd-7;
        fc1_weights[98][142] = 16'sd25;
        fc1_weights[98][143] = 16'sd1;
        fc1_weights[98][144] = 16'sd1;
        fc1_weights[98][145] = 16'sd27;
        fc1_weights[98][146] = 16'sd-7;
        fc1_weights[98][147] = 16'sd61;
        fc1_weights[98][148] = 16'sd11;
        fc1_weights[98][149] = 16'sd-17;
        fc1_weights[98][150] = 16'sd-1;
        fc1_weights[98][151] = 16'sd-10;
        fc1_weights[98][152] = 16'sd-29;
        fc1_weights[98][153] = 16'sd3;
        fc1_weights[98][154] = 16'sd-2;
        fc1_weights[98][155] = 16'sd-5;
        fc1_weights[98][156] = 16'sd24;
        fc1_weights[98][157] = 16'sd18;
        fc1_weights[98][158] = 16'sd12;
        fc1_weights[98][159] = 16'sd10;
        fc1_weights[98][160] = 16'sd-50;
        fc1_weights[98][161] = 16'sd-45;
        fc1_weights[98][162] = 16'sd-20;
        fc1_weights[98][163] = 16'sd-15;
        fc1_weights[98][164] = 16'sd-48;
        fc1_weights[98][165] = 16'sd-76;
        fc1_weights[98][166] = 16'sd-34;
        fc1_weights[98][167] = 16'sd3;
        fc1_weights[98][168] = 16'sd-46;
        fc1_weights[98][169] = 16'sd-1;
        fc1_weights[98][170] = 16'sd3;
        fc1_weights[98][171] = 16'sd-37;
        fc1_weights[98][172] = 16'sd-25;
        fc1_weights[98][173] = 16'sd-39;
        fc1_weights[98][174] = 16'sd-13;
        fc1_weights[98][175] = 16'sd-47;
        fc1_weights[98][176] = 16'sd-31;
        fc1_weights[98][177] = 16'sd-20;
        fc1_weights[98][178] = 16'sd-41;
        fc1_weights[98][179] = 16'sd-50;
        fc1_weights[98][180] = 16'sd-9;
        fc1_weights[98][181] = 16'sd13;
        fc1_weights[98][182] = 16'sd-34;
        fc1_weights[98][183] = 16'sd-1;
        fc1_weights[98][184] = 16'sd-43;
        fc1_weights[98][185] = 16'sd-48;
        fc1_weights[98][186] = 16'sd-37;
        fc1_weights[98][187] = 16'sd-18;
        fc1_weights[98][188] = 16'sd-56;
        fc1_weights[98][189] = 16'sd-39;
        fc1_weights[98][190] = 16'sd-26;
        fc1_weights[98][191] = 16'sd3;
        fc1_weights[98][192] = 16'sd-38;
        fc1_weights[98][193] = 16'sd-17;
        fc1_weights[98][194] = 16'sd-4;
        fc1_weights[98][195] = 16'sd18;
        fc1_weights[98][196] = 16'sd-5;
        fc1_weights[98][197] = 16'sd-28;
        fc1_weights[98][198] = 16'sd0;
        fc1_weights[98][199] = 16'sd1;
        fc1_weights[98][200] = 16'sd-8;
        fc1_weights[98][201] = 16'sd-30;
        fc1_weights[98][202] = 16'sd-33;
        fc1_weights[98][203] = 16'sd34;
        fc1_weights[98][204] = 16'sd-28;
        fc1_weights[98][205] = 16'sd14;
        fc1_weights[98][206] = 16'sd-12;
        fc1_weights[98][207] = 16'sd38;
        fc1_weights[99][0] = 16'sd14;
        fc1_weights[99][1] = 16'sd10;
        fc1_weights[99][2] = 16'sd-37;
        fc1_weights[99][3] = 16'sd-9;
        fc1_weights[99][4] = 16'sd-36;
        fc1_weights[99][5] = 16'sd8;
        fc1_weights[99][6] = 16'sd18;
        fc1_weights[99][7] = 16'sd-15;
        fc1_weights[99][8] = 16'sd-30;
        fc1_weights[99][9] = 16'sd-8;
        fc1_weights[99][10] = 16'sd33;
        fc1_weights[99][11] = 16'sd47;
        fc1_weights[99][12] = 16'sd83;
        fc1_weights[99][13] = 16'sd47;
        fc1_weights[99][14] = 16'sd100;
        fc1_weights[99][15] = 16'sd9;
        fc1_weights[99][16] = 16'sd-8;
        fc1_weights[99][17] = 16'sd-10;
        fc1_weights[99][18] = 16'sd-42;
        fc1_weights[99][19] = 16'sd1;
        fc1_weights[99][20] = 16'sd-97;
        fc1_weights[99][21] = 16'sd18;
        fc1_weights[99][22] = 16'sd39;
        fc1_weights[99][23] = 16'sd11;
        fc1_weights[99][24] = 16'sd-73;
        fc1_weights[99][25] = 16'sd-31;
        fc1_weights[99][26] = 16'sd-31;
        fc1_weights[99][27] = 16'sd-29;
        fc1_weights[99][28] = 16'sd-27;
        fc1_weights[99][29] = 16'sd-5;
        fc1_weights[99][30] = 16'sd-49;
        fc1_weights[99][31] = 16'sd-30;
        fc1_weights[99][32] = 16'sd-7;
        fc1_weights[99][33] = 16'sd22;
        fc1_weights[99][34] = 16'sd-4;
        fc1_weights[99][35] = 16'sd-20;
        fc1_weights[99][36] = 16'sd49;
        fc1_weights[99][37] = 16'sd121;
        fc1_weights[99][38] = 16'sd62;
        fc1_weights[99][39] = 16'sd19;
        fc1_weights[99][40] = 16'sd-18;
        fc1_weights[99][41] = 16'sd-70;
        fc1_weights[99][42] = 16'sd-51;
        fc1_weights[99][43] = 16'sd-45;
        fc1_weights[99][44] = 16'sd-34;
        fc1_weights[99][45] = 16'sd18;
        fc1_weights[99][46] = 16'sd-79;
        fc1_weights[99][47] = 16'sd-53;
        fc1_weights[99][48] = 16'sd-1;
        fc1_weights[99][49] = 16'sd-32;
        fc1_weights[99][50] = 16'sd49;
        fc1_weights[99][51] = 16'sd0;
        fc1_weights[99][52] = 16'sd42;
        fc1_weights[99][53] = 16'sd9;
        fc1_weights[99][54] = 16'sd44;
        fc1_weights[99][55] = 16'sd32;
        fc1_weights[99][56] = 16'sd37;
        fc1_weights[99][57] = 16'sd-31;
        fc1_weights[99][58] = 16'sd10;
        fc1_weights[99][59] = 16'sd-12;
        fc1_weights[99][60] = 16'sd34;
        fc1_weights[99][61] = 16'sd-48;
        fc1_weights[99][62] = 16'sd53;
        fc1_weights[99][63] = 16'sd39;
        fc1_weights[99][64] = 16'sd24;
        fc1_weights[99][65] = 16'sd-1;
        fc1_weights[99][66] = 16'sd-41;
        fc1_weights[99][67] = 16'sd-57;
        fc1_weights[99][68] = 16'sd-4;
        fc1_weights[99][69] = 16'sd57;
        fc1_weights[99][70] = 16'sd-4;
        fc1_weights[99][71] = 16'sd-104;
        fc1_weights[99][72] = 16'sd-84;
        fc1_weights[99][73] = 16'sd-6;
        fc1_weights[99][74] = 16'sd-5;
        fc1_weights[99][75] = 16'sd6;
        fc1_weights[99][76] = 16'sd8;
        fc1_weights[99][77] = 16'sd20;
        fc1_weights[99][78] = 16'sd4;
        fc1_weights[99][79] = 16'sd-19;
        fc1_weights[99][80] = 16'sd8;
        fc1_weights[99][81] = 16'sd24;
        fc1_weights[99][82] = 16'sd40;
        fc1_weights[99][83] = 16'sd37;
        fc1_weights[99][84] = 16'sd36;
        fc1_weights[99][85] = 16'sd17;
        fc1_weights[99][86] = 16'sd17;
        fc1_weights[99][87] = 16'sd-16;
        fc1_weights[99][88] = 16'sd-5;
        fc1_weights[99][89] = 16'sd-10;
        fc1_weights[99][90] = 16'sd-56;
        fc1_weights[99][91] = 16'sd-18;
        fc1_weights[99][92] = 16'sd-3;
        fc1_weights[99][93] = 16'sd-10;
        fc1_weights[99][94] = 16'sd76;
        fc1_weights[99][95] = 16'sd-3;
        fc1_weights[99][96] = 16'sd17;
        fc1_weights[99][97] = 16'sd-6;
        fc1_weights[99][98] = 16'sd-44;
        fc1_weights[99][99] = 16'sd7;
        fc1_weights[99][100] = 16'sd-8;
        fc1_weights[99][101] = 16'sd27;
        fc1_weights[99][102] = 16'sd16;
        fc1_weights[99][103] = 16'sd31;
        fc1_weights[99][104] = 16'sd2;
        fc1_weights[99][105] = 16'sd52;
        fc1_weights[99][106] = 16'sd33;
        fc1_weights[99][107] = 16'sd-17;
        fc1_weights[99][108] = 16'sd-45;
        fc1_weights[99][109] = 16'sd11;
        fc1_weights[99][110] = 16'sd-30;
        fc1_weights[99][111] = 16'sd12;
        fc1_weights[99][112] = 16'sd-37;
        fc1_weights[99][113] = 16'sd-25;
        fc1_weights[99][114] = 16'sd43;
        fc1_weights[99][115] = 16'sd67;
        fc1_weights[99][116] = 16'sd-22;
        fc1_weights[99][117] = 16'sd-92;
        fc1_weights[99][118] = 16'sd-45;
        fc1_weights[99][119] = 16'sd-39;
        fc1_weights[99][120] = 16'sd8;
        fc1_weights[99][121] = 16'sd-5;
        fc1_weights[99][122] = 16'sd-18;
        fc1_weights[99][123] = 16'sd-42;
        fc1_weights[99][124] = 16'sd1;
        fc1_weights[99][125] = 16'sd-10;
        fc1_weights[99][126] = 16'sd-12;
        fc1_weights[99][127] = 16'sd14;
        fc1_weights[99][128] = 16'sd13;
        fc1_weights[99][129] = 16'sd53;
        fc1_weights[99][130] = 16'sd22;
        fc1_weights[99][131] = 16'sd59;
        fc1_weights[99][132] = 16'sd-33;
        fc1_weights[99][133] = 16'sd-14;
        fc1_weights[99][134] = 16'sd-54;
        fc1_weights[99][135] = 16'sd2;
        fc1_weights[99][136] = 16'sd-4;
        fc1_weights[99][137] = 16'sd5;
        fc1_weights[99][138] = 16'sd21;
        fc1_weights[99][139] = 16'sd9;
        fc1_weights[99][140] = 16'sd-1;
        fc1_weights[99][141] = 16'sd39;
        fc1_weights[99][142] = 16'sd-48;
        fc1_weights[99][143] = 16'sd-4;
        fc1_weights[99][144] = 16'sd-45;
        fc1_weights[99][145] = 16'sd-62;
        fc1_weights[99][146] = 16'sd-32;
        fc1_weights[99][147] = 16'sd-61;
        fc1_weights[99][148] = 16'sd-79;
        fc1_weights[99][149] = 16'sd-61;
        fc1_weights[99][150] = 16'sd-22;
        fc1_weights[99][151] = 16'sd-28;
        fc1_weights[99][152] = 16'sd-1;
        fc1_weights[99][153] = 16'sd-1;
        fc1_weights[99][154] = 16'sd2;
        fc1_weights[99][155] = 16'sd-17;
        fc1_weights[99][156] = 16'sd-19;
        fc1_weights[99][157] = 16'sd4;
        fc1_weights[99][158] = 16'sd8;
        fc1_weights[99][159] = 16'sd-3;
        fc1_weights[99][160] = 16'sd68;
        fc1_weights[99][161] = 16'sd69;
        fc1_weights[99][162] = 16'sd16;
        fc1_weights[99][163] = 16'sd-4;
        fc1_weights[99][164] = 16'sd-17;
        fc1_weights[99][165] = 16'sd19;
        fc1_weights[99][166] = 16'sd10;
        fc1_weights[99][167] = 16'sd-14;
        fc1_weights[99][168] = 16'sd-19;
        fc1_weights[99][169] = 16'sd-28;
        fc1_weights[99][170] = 16'sd-62;
        fc1_weights[99][171] = 16'sd-13;
        fc1_weights[99][172] = 16'sd5;
        fc1_weights[99][173] = 16'sd-31;
        fc1_weights[99][174] = 16'sd30;
        fc1_weights[99][175] = 16'sd4;
        fc1_weights[99][176] = 16'sd18;
        fc1_weights[99][177] = 16'sd-17;
        fc1_weights[99][178] = 16'sd3;
        fc1_weights[99][179] = 16'sd35;
        fc1_weights[99][180] = 16'sd-14;
        fc1_weights[99][181] = 16'sd35;
        fc1_weights[99][182] = 16'sd69;
        fc1_weights[99][183] = 16'sd15;
        fc1_weights[99][184] = 16'sd14;
        fc1_weights[99][185] = 16'sd-36;
        fc1_weights[99][186] = 16'sd26;
        fc1_weights[99][187] = 16'sd20;
        fc1_weights[99][188] = 16'sd27;
        fc1_weights[99][189] = 16'sd-20;
        fc1_weights[99][190] = 16'sd-31;
        fc1_weights[99][191] = 16'sd-37;
        fc1_weights[99][192] = 16'sd29;
        fc1_weights[99][193] = 16'sd21;
        fc1_weights[99][194] = 16'sd-37;
        fc1_weights[99][195] = 16'sd-16;
        fc1_weights[99][196] = 16'sd-39;
        fc1_weights[99][197] = 16'sd-49;
        fc1_weights[99][198] = 16'sd-14;
        fc1_weights[99][199] = 16'sd-25;
        fc1_weights[99][200] = 16'sd6;
        fc1_weights[99][201] = 16'sd-7;
        fc1_weights[99][202] = 16'sd5;
        fc1_weights[99][203] = 16'sd52;
        fc1_weights[99][204] = 16'sd13;
        fc1_weights[99][205] = 16'sd-4;
        fc1_weights[99][206] = 16'sd32;
        fc1_weights[99][207] = 16'sd1;
        fc1_weights[100][0] = 16'sd-44;
        fc1_weights[100][1] = 16'sd47;
        fc1_weights[100][2] = 16'sd-23;
        fc1_weights[100][3] = 16'sd-27;
        fc1_weights[100][4] = 16'sd-80;
        fc1_weights[100][5] = 16'sd2;
        fc1_weights[100][6] = 16'sd-49;
        fc1_weights[100][7] = 16'sd66;
        fc1_weights[100][8] = 16'sd-49;
        fc1_weights[100][9] = 16'sd36;
        fc1_weights[100][10] = 16'sd91;
        fc1_weights[100][11] = 16'sd33;
        fc1_weights[100][12] = 16'sd-5;
        fc1_weights[100][13] = 16'sd-55;
        fc1_weights[100][14] = 16'sd-25;
        fc1_weights[100][15] = 16'sd11;
        fc1_weights[100][16] = 16'sd15;
        fc1_weights[100][17] = 16'sd9;
        fc1_weights[100][18] = 16'sd-2;
        fc1_weights[100][19] = 16'sd10;
        fc1_weights[100][20] = 16'sd67;
        fc1_weights[100][21] = 16'sd19;
        fc1_weights[100][22] = 16'sd-8;
        fc1_weights[100][23] = 16'sd-26;
        fc1_weights[100][24] = 16'sd13;
        fc1_weights[100][25] = 16'sd-17;
        fc1_weights[100][26] = 16'sd-16;
        fc1_weights[100][27] = 16'sd-24;
        fc1_weights[100][28] = 16'sd-36;
        fc1_weights[100][29] = 16'sd52;
        fc1_weights[100][30] = 16'sd-21;
        fc1_weights[100][31] = 16'sd9;
        fc1_weights[100][32] = 16'sd2;
        fc1_weights[100][33] = 16'sd-76;
        fc1_weights[100][34] = 16'sd10;
        fc1_weights[100][35] = 16'sd19;
        fc1_weights[100][36] = 16'sd75;
        fc1_weights[100][37] = 16'sd98;
        fc1_weights[100][38] = 16'sd53;
        fc1_weights[100][39] = 16'sd-79;
        fc1_weights[100][40] = 16'sd81;
        fc1_weights[100][41] = 16'sd-47;
        fc1_weights[100][42] = 16'sd15;
        fc1_weights[100][43] = 16'sd22;
        fc1_weights[100][44] = 16'sd29;
        fc1_weights[100][45] = 16'sd0;
        fc1_weights[100][46] = 16'sd-10;
        fc1_weights[100][47] = 16'sd9;
        fc1_weights[100][48] = 16'sd46;
        fc1_weights[100][49] = 16'sd59;
        fc1_weights[100][50] = 16'sd-30;
        fc1_weights[100][51] = 16'sd-77;
        fc1_weights[100][52] = 16'sd-37;
        fc1_weights[100][53] = 16'sd-10;
        fc1_weights[100][54] = 16'sd39;
        fc1_weights[100][55] = 16'sd18;
        fc1_weights[100][56] = 16'sd29;
        fc1_weights[100][57] = 16'sd63;
        fc1_weights[100][58] = 16'sd-7;
        fc1_weights[100][59] = 16'sd-62;
        fc1_weights[100][60] = 16'sd66;
        fc1_weights[100][61] = 16'sd69;
        fc1_weights[100][62] = 16'sd-4;
        fc1_weights[100][63] = 16'sd42;
        fc1_weights[100][64] = 16'sd121;
        fc1_weights[100][65] = 16'sd-109;
        fc1_weights[100][66] = 16'sd1;
        fc1_weights[100][67] = 16'sd-63;
        fc1_weights[100][68] = 16'sd-16;
        fc1_weights[100][69] = 16'sd57;
        fc1_weights[100][70] = 16'sd-4;
        fc1_weights[100][71] = 16'sd28;
        fc1_weights[100][72] = 16'sd39;
        fc1_weights[100][73] = 16'sd3;
        fc1_weights[100][74] = 16'sd15;
        fc1_weights[100][75] = 16'sd-30;
        fc1_weights[100][76] = 16'sd17;
        fc1_weights[100][77] = 16'sd30;
        fc1_weights[100][78] = 16'sd-14;
        fc1_weights[100][79] = 16'sd35;
        fc1_weights[100][80] = 16'sd13;
        fc1_weights[100][81] = 16'sd-13;
        fc1_weights[100][82] = 16'sd-35;
        fc1_weights[100][83] = 16'sd-18;
        fc1_weights[100][84] = 16'sd11;
        fc1_weights[100][85] = 16'sd-72;
        fc1_weights[100][86] = 16'sd-4;
        fc1_weights[100][87] = 16'sd65;
        fc1_weights[100][88] = 16'sd1;
        fc1_weights[100][89] = 16'sd-3;
        fc1_weights[100][90] = 16'sd11;
        fc1_weights[100][91] = 16'sd31;
        fc1_weights[100][92] = 16'sd14;
        fc1_weights[100][93] = 16'sd-10;
        fc1_weights[100][94] = 16'sd18;
        fc1_weights[100][95] = 16'sd51;
        fc1_weights[100][96] = 16'sd-7;
        fc1_weights[100][97] = 16'sd-10;
        fc1_weights[100][98] = 16'sd26;
        fc1_weights[100][99] = 16'sd-38;
        fc1_weights[100][100] = 16'sd-2;
        fc1_weights[100][101] = 16'sd20;
        fc1_weights[100][102] = 16'sd-21;
        fc1_weights[100][103] = 16'sd-29;
        fc1_weights[100][104] = 16'sd-6;
        fc1_weights[100][105] = 16'sd-19;
        fc1_weights[100][106] = 16'sd8;
        fc1_weights[100][107] = 16'sd-42;
        fc1_weights[100][108] = 16'sd-44;
        fc1_weights[100][109] = 16'sd-68;
        fc1_weights[100][110] = 16'sd-28;
        fc1_weights[100][111] = 16'sd-20;
        fc1_weights[100][112] = 16'sd21;
        fc1_weights[100][113] = 16'sd-5;
        fc1_weights[100][114] = 16'sd54;
        fc1_weights[100][115] = 16'sd31;
        fc1_weights[100][116] = 16'sd34;
        fc1_weights[100][117] = 16'sd94;
        fc1_weights[100][118] = 16'sd68;
        fc1_weights[100][119] = 16'sd5;
        fc1_weights[100][120] = 16'sd-44;
        fc1_weights[100][121] = 16'sd94;
        fc1_weights[100][122] = 16'sd8;
        fc1_weights[100][123] = 16'sd-58;
        fc1_weights[100][124] = 16'sd-53;
        fc1_weights[100][125] = 16'sd-9;
        fc1_weights[100][126] = 16'sd-28;
        fc1_weights[100][127] = 16'sd28;
        fc1_weights[100][128] = 16'sd-38;
        fc1_weights[100][129] = 16'sd-94;
        fc1_weights[100][130] = 16'sd-52;
        fc1_weights[100][131] = 16'sd-11;
        fc1_weights[100][132] = 16'sd4;
        fc1_weights[100][133] = 16'sd-50;
        fc1_weights[100][134] = 16'sd-10;
        fc1_weights[100][135] = 16'sd16;
        fc1_weights[100][136] = 16'sd-11;
        fc1_weights[100][137] = 16'sd-26;
        fc1_weights[100][138] = 16'sd100;
        fc1_weights[100][139] = 16'sd-30;
        fc1_weights[100][140] = 16'sd-56;
        fc1_weights[100][141] = 16'sd-50;
        fc1_weights[100][142] = 16'sd46;
        fc1_weights[100][143] = 16'sd27;
        fc1_weights[100][144] = 16'sd63;
        fc1_weights[100][145] = 16'sd15;
        fc1_weights[100][146] = 16'sd32;
        fc1_weights[100][147] = 16'sd43;
        fc1_weights[100][148] = 16'sd-35;
        fc1_weights[100][149] = 16'sd9;
        fc1_weights[100][150] = 16'sd-23;
        fc1_weights[100][151] = 16'sd1;
        fc1_weights[100][152] = 16'sd34;
        fc1_weights[100][153] = 16'sd17;
        fc1_weights[100][154] = 16'sd-35;
        fc1_weights[100][155] = 16'sd5;
        fc1_weights[100][156] = 16'sd-53;
        fc1_weights[100][157] = 16'sd9;
        fc1_weights[100][158] = 16'sd-39;
        fc1_weights[100][159] = 16'sd12;
        fc1_weights[100][160] = 16'sd-57;
        fc1_weights[100][161] = 16'sd-49;
        fc1_weights[100][162] = 16'sd47;
        fc1_weights[100][163] = 16'sd-45;
        fc1_weights[100][164] = 16'sd-63;
        fc1_weights[100][165] = 16'sd-15;
        fc1_weights[100][166] = 16'sd9;
        fc1_weights[100][167] = 16'sd-9;
        fc1_weights[100][168] = 16'sd39;
        fc1_weights[100][169] = 16'sd-4;
        fc1_weights[100][170] = 16'sd11;
        fc1_weights[100][171] = 16'sd-65;
        fc1_weights[100][172] = 16'sd42;
        fc1_weights[100][173] = 16'sd-18;
        fc1_weights[100][174] = 16'sd0;
        fc1_weights[100][175] = 16'sd-6;
        fc1_weights[100][176] = 16'sd-37;
        fc1_weights[100][177] = 16'sd16;
        fc1_weights[100][178] = 16'sd-33;
        fc1_weights[100][179] = 16'sd51;
        fc1_weights[100][180] = 16'sd4;
        fc1_weights[100][181] = 16'sd10;
        fc1_weights[100][182] = 16'sd11;
        fc1_weights[100][183] = 16'sd-30;
        fc1_weights[100][184] = 16'sd-12;
        fc1_weights[100][185] = 16'sd61;
        fc1_weights[100][186] = 16'sd-34;
        fc1_weights[100][187] = 16'sd-7;
        fc1_weights[100][188] = 16'sd1;
        fc1_weights[100][189] = 16'sd-74;
        fc1_weights[100][190] = 16'sd6;
        fc1_weights[100][191] = 16'sd76;
        fc1_weights[100][192] = 16'sd-20;
        fc1_weights[100][193] = 16'sd-38;
        fc1_weights[100][194] = 16'sd-51;
        fc1_weights[100][195] = 16'sd-7;
        fc1_weights[100][196] = 16'sd-41;
        fc1_weights[100][197] = 16'sd56;
        fc1_weights[100][198] = 16'sd-19;
        fc1_weights[100][199] = 16'sd-30;
        fc1_weights[100][200] = 16'sd37;
        fc1_weights[100][201] = 16'sd16;
        fc1_weights[100][202] = 16'sd-9;
        fc1_weights[100][203] = 16'sd21;
        fc1_weights[100][204] = 16'sd83;
        fc1_weights[100][205] = 16'sd43;
        fc1_weights[100][206] = 16'sd-9;
        fc1_weights[100][207] = 16'sd2;
        fc1_weights[101][0] = 16'sd58;
        fc1_weights[101][1] = 16'sd52;
        fc1_weights[101][2] = 16'sd14;
        fc1_weights[101][3] = 16'sd25;
        fc1_weights[101][4] = 16'sd-1;
        fc1_weights[101][5] = 16'sd-2;
        fc1_weights[101][6] = 16'sd36;
        fc1_weights[101][7] = 16'sd29;
        fc1_weights[101][8] = 16'sd-17;
        fc1_weights[101][9] = 16'sd-7;
        fc1_weights[101][10] = 16'sd7;
        fc1_weights[101][11] = 16'sd-38;
        fc1_weights[101][12] = 16'sd-47;
        fc1_weights[101][13] = 16'sd-21;
        fc1_weights[101][14] = 16'sd-37;
        fc1_weights[101][15] = 16'sd-62;
        fc1_weights[101][16] = 16'sd-14;
        fc1_weights[101][17] = 16'sd-47;
        fc1_weights[101][18] = 16'sd-24;
        fc1_weights[101][19] = 16'sd-3;
        fc1_weights[101][20] = 16'sd17;
        fc1_weights[101][21] = 16'sd40;
        fc1_weights[101][22] = 16'sd33;
        fc1_weights[101][23] = 16'sd-1;
        fc1_weights[101][24] = 16'sd32;
        fc1_weights[101][25] = 16'sd14;
        fc1_weights[101][26] = 16'sd7;
        fc1_weights[101][27] = 16'sd8;
        fc1_weights[101][28] = 16'sd42;
        fc1_weights[101][29] = 16'sd22;
        fc1_weights[101][30] = 16'sd-30;
        fc1_weights[101][31] = 16'sd-9;
        fc1_weights[101][32] = 16'sd40;
        fc1_weights[101][33] = 16'sd54;
        fc1_weights[101][34] = 16'sd10;
        fc1_weights[101][35] = 16'sd2;
        fc1_weights[101][36] = 16'sd-3;
        fc1_weights[101][37] = 16'sd-28;
        fc1_weights[101][38] = 16'sd-57;
        fc1_weights[101][39] = 16'sd-38;
        fc1_weights[101][40] = 16'sd-60;
        fc1_weights[101][41] = 16'sd-7;
        fc1_weights[101][42] = 16'sd-35;
        fc1_weights[101][43] = 16'sd2;
        fc1_weights[101][44] = 16'sd0;
        fc1_weights[101][45] = 16'sd7;
        fc1_weights[101][46] = 16'sd18;
        fc1_weights[101][47] = 16'sd50;
        fc1_weights[101][48] = 16'sd9;
        fc1_weights[101][49] = 16'sd-23;
        fc1_weights[101][50] = 16'sd18;
        fc1_weights[101][51] = 16'sd25;
        fc1_weights[101][52] = 16'sd-52;
        fc1_weights[101][53] = 16'sd-19;
        fc1_weights[101][54] = 16'sd41;
        fc1_weights[101][55] = 16'sd36;
        fc1_weights[101][56] = 16'sd-12;
        fc1_weights[101][57] = 16'sd23;
        fc1_weights[101][58] = 16'sd45;
        fc1_weights[101][59] = 16'sd22;
        fc1_weights[101][60] = 16'sd-7;
        fc1_weights[101][61] = 16'sd20;
        fc1_weights[101][62] = 16'sd15;
        fc1_weights[101][63] = 16'sd-45;
        fc1_weights[101][64] = 16'sd-39;
        fc1_weights[101][65] = 16'sd-5;
        fc1_weights[101][66] = 16'sd-16;
        fc1_weights[101][67] = 16'sd-12;
        fc1_weights[101][68] = 16'sd-11;
        fc1_weights[101][69] = 16'sd31;
        fc1_weights[101][70] = 16'sd-23;
        fc1_weights[101][71] = 16'sd-8;
        fc1_weights[101][72] = 16'sd39;
        fc1_weights[101][73] = 16'sd-13;
        fc1_weights[101][74] = 16'sd-13;
        fc1_weights[101][75] = 16'sd-46;
        fc1_weights[101][76] = 16'sd-10;
        fc1_weights[101][77] = 16'sd38;
        fc1_weights[101][78] = 16'sd-96;
        fc1_weights[101][79] = 16'sd-70;
        fc1_weights[101][80] = 16'sd-39;
        fc1_weights[101][81] = 16'sd11;
        fc1_weights[101][82] = 16'sd18;
        fc1_weights[101][83] = 16'sd-5;
        fc1_weights[101][84] = 16'sd41;
        fc1_weights[101][85] = 16'sd80;
        fc1_weights[101][86] = 16'sd-3;
        fc1_weights[101][87] = 16'sd-37;
        fc1_weights[101][88] = 16'sd24;
        fc1_weights[101][89] = 16'sd-13;
        fc1_weights[101][90] = 16'sd-41;
        fc1_weights[101][91] = 16'sd-20;
        fc1_weights[101][92] = 16'sd4;
        fc1_weights[101][93] = 16'sd19;
        fc1_weights[101][94] = 16'sd29;
        fc1_weights[101][95] = 16'sd10;
        fc1_weights[101][96] = 16'sd-13;
        fc1_weights[101][97] = 16'sd-16;
        fc1_weights[101][98] = 16'sd-21;
        fc1_weights[101][99] = 16'sd-13;
        fc1_weights[101][100] = 16'sd-13;
        fc1_weights[101][101] = 16'sd27;
        fc1_weights[101][102] = 16'sd68;
        fc1_weights[101][103] = 16'sd44;
        fc1_weights[101][104] = 16'sd-61;
        fc1_weights[101][105] = 16'sd-51;
        fc1_weights[101][106] = 16'sd-11;
        fc1_weights[101][107] = 16'sd-4;
        fc1_weights[101][108] = 16'sd-20;
        fc1_weights[101][109] = 16'sd-12;
        fc1_weights[101][110] = 16'sd-34;
        fc1_weights[101][111] = 16'sd2;
        fc1_weights[101][112] = 16'sd-33;
        fc1_weights[101][113] = 16'sd-58;
        fc1_weights[101][114] = 16'sd-1;
        fc1_weights[101][115] = 16'sd-12;
        fc1_weights[101][116] = 16'sd6;
        fc1_weights[101][117] = 16'sd-27;
        fc1_weights[101][118] = 16'sd-56;
        fc1_weights[101][119] = 16'sd-58;
        fc1_weights[101][120] = 16'sd-37;
        fc1_weights[101][121] = 16'sd-5;
        fc1_weights[101][122] = 16'sd11;
        fc1_weights[101][123] = 16'sd-43;
        fc1_weights[101][124] = 16'sd-38;
        fc1_weights[101][125] = 16'sd-14;
        fc1_weights[101][126] = 16'sd15;
        fc1_weights[101][127] = 16'sd-16;
        fc1_weights[101][128] = 16'sd-11;
        fc1_weights[101][129] = 16'sd27;
        fc1_weights[101][130] = 16'sd-44;
        fc1_weights[101][131] = 16'sd-46;
        fc1_weights[101][132] = 16'sd-27;
        fc1_weights[101][133] = 16'sd-73;
        fc1_weights[101][134] = 16'sd-20;
        fc1_weights[101][135] = 16'sd-22;
        fc1_weights[101][136] = 16'sd-27;
        fc1_weights[101][137] = 16'sd-47;
        fc1_weights[101][138] = 16'sd-50;
        fc1_weights[101][139] = 16'sd9;
        fc1_weights[101][140] = 16'sd39;
        fc1_weights[101][141] = 16'sd-16;
        fc1_weights[101][142] = 16'sd-33;
        fc1_weights[101][143] = 16'sd42;
        fc1_weights[101][144] = 16'sd-16;
        fc1_weights[101][145] = 16'sd8;
        fc1_weights[101][146] = 16'sd-19;
        fc1_weights[101][147] = 16'sd-19;
        fc1_weights[101][148] = 16'sd-35;
        fc1_weights[101][149] = 16'sd4;
        fc1_weights[101][150] = 16'sd4;
        fc1_weights[101][151] = 16'sd34;
        fc1_weights[101][152] = 16'sd25;
        fc1_weights[101][153] = 16'sd19;
        fc1_weights[101][154] = 16'sd-9;
        fc1_weights[101][155] = 16'sd54;
        fc1_weights[101][156] = 16'sd-5;
        fc1_weights[101][157] = 16'sd-28;
        fc1_weights[101][158] = 16'sd-16;
        fc1_weights[101][159] = 16'sd8;
        fc1_weights[101][160] = 16'sd-13;
        fc1_weights[101][161] = 16'sd-41;
        fc1_weights[101][162] = 16'sd-77;
        fc1_weights[101][163] = 16'sd-16;
        fc1_weights[101][164] = 16'sd21;
        fc1_weights[101][165] = 16'sd13;
        fc1_weights[101][166] = 16'sd11;
        fc1_weights[101][167] = 16'sd10;
        fc1_weights[101][168] = 16'sd-12;
        fc1_weights[101][169] = 16'sd-25;
        fc1_weights[101][170] = 16'sd-33;
        fc1_weights[101][171] = 16'sd-32;
        fc1_weights[101][172] = 16'sd-7;
        fc1_weights[101][173] = 16'sd-29;
        fc1_weights[101][174] = 16'sd-32;
        fc1_weights[101][175] = 16'sd-7;
        fc1_weights[101][176] = 16'sd33;
        fc1_weights[101][177] = 16'sd31;
        fc1_weights[101][178] = 16'sd50;
        fc1_weights[101][179] = 16'sd60;
        fc1_weights[101][180] = 16'sd35;
        fc1_weights[101][181] = 16'sd82;
        fc1_weights[101][182] = 16'sd-17;
        fc1_weights[101][183] = 16'sd10;
        fc1_weights[101][184] = 16'sd28;
        fc1_weights[101][185] = 16'sd-1;
        fc1_weights[101][186] = 16'sd-30;
        fc1_weights[101][187] = 16'sd-25;
        fc1_weights[101][188] = 16'sd19;
        fc1_weights[101][189] = 16'sd19;
        fc1_weights[101][190] = 16'sd-3;
        fc1_weights[101][191] = 16'sd35;
        fc1_weights[101][192] = 16'sd63;
        fc1_weights[101][193] = 16'sd51;
        fc1_weights[101][194] = 16'sd1;
        fc1_weights[101][195] = 16'sd32;
        fc1_weights[101][196] = 16'sd35;
        fc1_weights[101][197] = 16'sd6;
        fc1_weights[101][198] = 16'sd63;
        fc1_weights[101][199] = 16'sd37;
        fc1_weights[101][200] = 16'sd34;
        fc1_weights[101][201] = 16'sd45;
        fc1_weights[101][202] = 16'sd1;
        fc1_weights[101][203] = 16'sd31;
        fc1_weights[101][204] = 16'sd64;
        fc1_weights[101][205] = 16'sd82;
        fc1_weights[101][206] = 16'sd66;
        fc1_weights[101][207] = 16'sd64;
        fc1_weights[102][0] = 16'sd9;
        fc1_weights[102][1] = 16'sd53;
        fc1_weights[102][2] = 16'sd-20;
        fc1_weights[102][3] = 16'sd-11;
        fc1_weights[102][4] = 16'sd-31;
        fc1_weights[102][5] = 16'sd-28;
        fc1_weights[102][6] = 16'sd-84;
        fc1_weights[102][7] = 16'sd25;
        fc1_weights[102][8] = 16'sd-69;
        fc1_weights[102][9] = 16'sd-16;
        fc1_weights[102][10] = 16'sd-2;
        fc1_weights[102][11] = 16'sd-80;
        fc1_weights[102][12] = 16'sd-89;
        fc1_weights[102][13] = 16'sd-5;
        fc1_weights[102][14] = 16'sd35;
        fc1_weights[102][15] = 16'sd59;
        fc1_weights[102][16] = 16'sd-7;
        fc1_weights[102][17] = 16'sd-30;
        fc1_weights[102][18] = 16'sd1;
        fc1_weights[102][19] = 16'sd40;
        fc1_weights[102][20] = 16'sd49;
        fc1_weights[102][21] = 16'sd91;
        fc1_weights[102][22] = 16'sd58;
        fc1_weights[102][23] = 16'sd1;
        fc1_weights[102][24] = 16'sd21;
        fc1_weights[102][25] = 16'sd29;
        fc1_weights[102][26] = 16'sd21;
        fc1_weights[102][27] = 16'sd29;
        fc1_weights[102][28] = 16'sd25;
        fc1_weights[102][29] = 16'sd45;
        fc1_weights[102][30] = 16'sd23;
        fc1_weights[102][31] = 16'sd-66;
        fc1_weights[102][32] = 16'sd-63;
        fc1_weights[102][33] = 16'sd-80;
        fc1_weights[102][34] = 16'sd-76;
        fc1_weights[102][35] = 16'sd-36;
        fc1_weights[102][36] = 16'sd22;
        fc1_weights[102][37] = 16'sd31;
        fc1_weights[102][38] = 16'sd-2;
        fc1_weights[102][39] = 16'sd38;
        fc1_weights[102][40] = 16'sd97;
        fc1_weights[102][41] = 16'sd4;
        fc1_weights[102][42] = 16'sd-95;
        fc1_weights[102][43] = 16'sd-7;
        fc1_weights[102][44] = 16'sd-3;
        fc1_weights[102][45] = 16'sd-7;
        fc1_weights[102][46] = 16'sd-80;
        fc1_weights[102][47] = 16'sd4;
        fc1_weights[102][48] = 16'sd77;
        fc1_weights[102][49] = 16'sd32;
        fc1_weights[102][50] = 16'sd36;
        fc1_weights[102][51] = 16'sd-93;
        fc1_weights[102][52] = 16'sd8;
        fc1_weights[102][53] = 16'sd24;
        fc1_weights[102][54] = 16'sd9;
        fc1_weights[102][55] = 16'sd47;
        fc1_weights[102][56] = 16'sd12;
        fc1_weights[102][57] = 16'sd-16;
        fc1_weights[102][58] = 16'sd-3;
        fc1_weights[102][59] = 16'sd-18;
        fc1_weights[102][60] = 16'sd-23;
        fc1_weights[102][61] = 16'sd27;
        fc1_weights[102][62] = 16'sd-104;
        fc1_weights[102][63] = 16'sd-45;
        fc1_weights[102][64] = 16'sd41;
        fc1_weights[102][65] = 16'sd-85;
        fc1_weights[102][66] = 16'sd-11;
        fc1_weights[102][67] = 16'sd8;
        fc1_weights[102][68] = 16'sd-118;
        fc1_weights[102][69] = 16'sd46;
        fc1_weights[102][70] = 16'sd4;
        fc1_weights[102][71] = 16'sd86;
        fc1_weights[102][72] = 16'sd34;
        fc1_weights[102][73] = 16'sd-29;
        fc1_weights[102][74] = 16'sd-19;
        fc1_weights[102][75] = 16'sd12;
        fc1_weights[102][76] = 16'sd-25;
        fc1_weights[102][77] = 16'sd-26;
        fc1_weights[102][78] = 16'sd23;
        fc1_weights[102][79] = 16'sd54;
        fc1_weights[102][80] = 16'sd46;
        fc1_weights[102][81] = 16'sd31;
        fc1_weights[102][82] = 16'sd24;
        fc1_weights[102][83] = 16'sd-54;
        fc1_weights[102][84] = 16'sd5;
        fc1_weights[102][85] = 16'sd-16;
        fc1_weights[102][86] = 16'sd-32;
        fc1_weights[102][87] = 16'sd27;
        fc1_weights[102][88] = 16'sd27;
        fc1_weights[102][89] = 16'sd41;
        fc1_weights[102][90] = 16'sd114;
        fc1_weights[102][91] = 16'sd126;
        fc1_weights[102][92] = 16'sd81;
        fc1_weights[102][93] = 16'sd57;
        fc1_weights[102][94] = 16'sd-75;
        fc1_weights[102][95] = 16'sd-49;
        fc1_weights[102][96] = 16'sd-13;
        fc1_weights[102][97] = 16'sd10;
        fc1_weights[102][98] = 16'sd19;
        fc1_weights[102][99] = 16'sd-10;
        fc1_weights[102][100] = 16'sd40;
        fc1_weights[102][101] = 16'sd19;
        fc1_weights[102][102] = 16'sd-57;
        fc1_weights[102][103] = 16'sd-112;
        fc1_weights[102][104] = 16'sd74;
        fc1_weights[102][105] = 16'sd-44;
        fc1_weights[102][106] = 16'sd0;
        fc1_weights[102][107] = 16'sd6;
        fc1_weights[102][108] = 16'sd-20;
        fc1_weights[102][109] = 16'sd1;
        fc1_weights[102][110] = 16'sd62;
        fc1_weights[102][111] = 16'sd32;
        fc1_weights[102][112] = 16'sd8;
        fc1_weights[102][113] = 16'sd-33;
        fc1_weights[102][114] = 16'sd-47;
        fc1_weights[102][115] = 16'sd-27;
        fc1_weights[102][116] = 16'sd-28;
        fc1_weights[102][117] = 16'sd16;
        fc1_weights[102][118] = 16'sd24;
        fc1_weights[102][119] = 16'sd-44;
        fc1_weights[102][120] = 16'sd-86;
        fc1_weights[102][121] = 16'sd-56;
        fc1_weights[102][122] = 16'sd27;
        fc1_weights[102][123] = 16'sd25;
        fc1_weights[102][124] = 16'sd-94;
        fc1_weights[102][125] = 16'sd-44;
        fc1_weights[102][126] = 16'sd-53;
        fc1_weights[102][127] = 16'sd10;
        fc1_weights[102][128] = 16'sd-78;
        fc1_weights[102][129] = 16'sd-128;
        fc1_weights[102][130] = 16'sd6;
        fc1_weights[102][131] = 16'sd-40;
        fc1_weights[102][132] = 16'sd-4;
        fc1_weights[102][133] = 16'sd33;
        fc1_weights[102][134] = 16'sd39;
        fc1_weights[102][135] = 16'sd9;
        fc1_weights[102][136] = 16'sd112;
        fc1_weights[102][137] = 16'sd105;
        fc1_weights[102][138] = 16'sd58;
        fc1_weights[102][139] = 16'sd-37;
        fc1_weights[102][140] = 16'sd-19;
        fc1_weights[102][141] = 16'sd-19;
        fc1_weights[102][142] = 16'sd34;
        fc1_weights[102][143] = 16'sd-15;
        fc1_weights[102][144] = 16'sd-46;
        fc1_weights[102][145] = 16'sd-8;
        fc1_weights[102][146] = 16'sd-24;
        fc1_weights[102][147] = 16'sd42;
        fc1_weights[102][148] = 16'sd37;
        fc1_weights[102][149] = 16'sd-38;
        fc1_weights[102][150] = 16'sd-20;
        fc1_weights[102][151] = 16'sd-28;
        fc1_weights[102][152] = 16'sd-18;
        fc1_weights[102][153] = 16'sd33;
        fc1_weights[102][154] = 16'sd-13;
        fc1_weights[102][155] = 16'sd6;
        fc1_weights[102][156] = 16'sd25;
        fc1_weights[102][157] = 16'sd55;
        fc1_weights[102][158] = 16'sd4;
        fc1_weights[102][159] = 16'sd-6;
        fc1_weights[102][160] = 16'sd33;
        fc1_weights[102][161] = 16'sd8;
        fc1_weights[102][162] = 16'sd38;
        fc1_weights[102][163] = 16'sd-15;
        fc1_weights[102][164] = 16'sd4;
        fc1_weights[102][165] = 16'sd-87;
        fc1_weights[102][166] = 16'sd-2;
        fc1_weights[102][167] = 16'sd32;
        fc1_weights[102][168] = 16'sd-27;
        fc1_weights[102][169] = 16'sd-5;
        fc1_weights[102][170] = 16'sd-31;
        fc1_weights[102][171] = 16'sd10;
        fc1_weights[102][172] = 16'sd53;
        fc1_weights[102][173] = 16'sd13;
        fc1_weights[102][174] = 16'sd-24;
        fc1_weights[102][175] = 16'sd-34;
        fc1_weights[102][176] = 16'sd-45;
        fc1_weights[102][177] = 16'sd-20;
        fc1_weights[102][178] = 16'sd-60;
        fc1_weights[102][179] = 16'sd-18;
        fc1_weights[102][180] = 16'sd-36;
        fc1_weights[102][181] = 16'sd-23;
        fc1_weights[102][182] = 16'sd25;
        fc1_weights[102][183] = 16'sd27;
        fc1_weights[102][184] = 16'sd-19;
        fc1_weights[102][185] = 16'sd47;
        fc1_weights[102][186] = 16'sd45;
        fc1_weights[102][187] = 16'sd47;
        fc1_weights[102][188] = 16'sd-56;
        fc1_weights[102][189] = 16'sd-7;
        fc1_weights[102][190] = 16'sd-21;
        fc1_weights[102][191] = 16'sd24;
        fc1_weights[102][192] = 16'sd-65;
        fc1_weights[102][193] = 16'sd-5;
        fc1_weights[102][194] = 16'sd9;
        fc1_weights[102][195] = 16'sd-9;
        fc1_weights[102][196] = 16'sd-31;
        fc1_weights[102][197] = 16'sd31;
        fc1_weights[102][198] = 16'sd-29;
        fc1_weights[102][199] = 16'sd25;
        fc1_weights[102][200] = 16'sd41;
        fc1_weights[102][201] = 16'sd-4;
        fc1_weights[102][202] = 16'sd52;
        fc1_weights[102][203] = 16'sd43;
        fc1_weights[102][204] = 16'sd33;
        fc1_weights[102][205] = 16'sd23;
        fc1_weights[102][206] = 16'sd-26;
        fc1_weights[102][207] = 16'sd-27;
        fc1_weights[103][0] = 16'sd22;
        fc1_weights[103][1] = 16'sd-2;
        fc1_weights[103][2] = 16'sd-11;
        fc1_weights[103][3] = 16'sd9;
        fc1_weights[103][4] = 16'sd16;
        fc1_weights[103][5] = 16'sd29;
        fc1_weights[103][6] = 16'sd32;
        fc1_weights[103][7] = 16'sd-45;
        fc1_weights[103][8] = 16'sd1;
        fc1_weights[103][9] = 16'sd-32;
        fc1_weights[103][10] = 16'sd-61;
        fc1_weights[103][11] = 16'sd-8;
        fc1_weights[103][12] = 16'sd-19;
        fc1_weights[103][13] = 16'sd-29;
        fc1_weights[103][14] = 16'sd-19;
        fc1_weights[103][15] = 16'sd18;
        fc1_weights[103][16] = 16'sd-18;
        fc1_weights[103][17] = 16'sd-39;
        fc1_weights[103][18] = 16'sd25;
        fc1_weights[103][19] = 16'sd-18;
        fc1_weights[103][20] = 16'sd22;
        fc1_weights[103][21] = 16'sd10;
        fc1_weights[103][22] = 16'sd3;
        fc1_weights[103][23] = 16'sd42;
        fc1_weights[103][24] = 16'sd100;
        fc1_weights[103][25] = 16'sd34;
        fc1_weights[103][26] = 16'sd5;
        fc1_weights[103][27] = 16'sd-9;
        fc1_weights[103][28] = 16'sd15;
        fc1_weights[103][29] = 16'sd36;
        fc1_weights[103][30] = 16'sd39;
        fc1_weights[103][31] = 16'sd61;
        fc1_weights[103][32] = 16'sd24;
        fc1_weights[103][33] = 16'sd-48;
        fc1_weights[103][34] = 16'sd0;
        fc1_weights[103][35] = 16'sd1;
        fc1_weights[103][36] = 16'sd25;
        fc1_weights[103][37] = 16'sd7;
        fc1_weights[103][38] = 16'sd-23;
        fc1_weights[103][39] = 16'sd-3;
        fc1_weights[103][40] = 16'sd3;
        fc1_weights[103][41] = 16'sd-23;
        fc1_weights[103][42] = 16'sd33;
        fc1_weights[103][43] = 16'sd-47;
        fc1_weights[103][44] = 16'sd-5;
        fc1_weights[103][45] = 16'sd0;
        fc1_weights[103][46] = 16'sd-34;
        fc1_weights[103][47] = 16'sd-37;
        fc1_weights[103][48] = 16'sd-26;
        fc1_weights[103][49] = 16'sd56;
        fc1_weights[103][50] = 16'sd26;
        fc1_weights[103][51] = 16'sd9;
        fc1_weights[103][52] = 16'sd18;
        fc1_weights[103][53] = 16'sd-29;
        fc1_weights[103][54] = 16'sd18;
        fc1_weights[103][55] = 16'sd-1;
        fc1_weights[103][56] = 16'sd9;
        fc1_weights[103][57] = 16'sd-1;
        fc1_weights[103][58] = 16'sd19;
        fc1_weights[103][59] = 16'sd60;
        fc1_weights[103][60] = 16'sd78;
        fc1_weights[103][61] = 16'sd-7;
        fc1_weights[103][62] = 16'sd-7;
        fc1_weights[103][63] = 16'sd-15;
        fc1_weights[103][64] = 16'sd36;
        fc1_weights[103][65] = 16'sd26;
        fc1_weights[103][66] = 16'sd-27;
        fc1_weights[103][67] = 16'sd-67;
        fc1_weights[103][68] = 16'sd-67;
        fc1_weights[103][69] = 16'sd-65;
        fc1_weights[103][70] = 16'sd-5;
        fc1_weights[103][71] = 16'sd36;
        fc1_weights[103][72] = 16'sd-9;
        fc1_weights[103][73] = 16'sd-36;
        fc1_weights[103][74] = 16'sd-52;
        fc1_weights[103][75] = 16'sd-17;
        fc1_weights[103][76] = 16'sd18;
        fc1_weights[103][77] = 16'sd16;
        fc1_weights[103][78] = 16'sd63;
        fc1_weights[103][79] = 16'sd55;
        fc1_weights[103][80] = 16'sd0;
        fc1_weights[103][81] = 16'sd-49;
        fc1_weights[103][82] = 16'sd-1;
        fc1_weights[103][83] = 16'sd24;
        fc1_weights[103][84] = 16'sd18;
        fc1_weights[103][85] = 16'sd-20;
        fc1_weights[103][86] = 16'sd13;
        fc1_weights[103][87] = 16'sd36;
        fc1_weights[103][88] = 16'sd-39;
        fc1_weights[103][89] = 16'sd18;
        fc1_weights[103][90] = 16'sd100;
        fc1_weights[103][91] = 16'sd-26;
        fc1_weights[103][92] = 16'sd-5;
        fc1_weights[103][93] = 16'sd-34;
        fc1_weights[103][94] = 16'sd-79;
        fc1_weights[103][95] = 16'sd-41;
        fc1_weights[103][96] = 16'sd-5;
        fc1_weights[103][97] = 16'sd-23;
        fc1_weights[103][98] = 16'sd-30;
        fc1_weights[103][99] = 16'sd-37;
        fc1_weights[103][100] = 16'sd1;
        fc1_weights[103][101] = 16'sd8;
        fc1_weights[103][102] = 16'sd-25;
        fc1_weights[103][103] = 16'sd-45;
        fc1_weights[103][104] = 16'sd46;
        fc1_weights[103][105] = 16'sd10;
        fc1_weights[103][106] = 16'sd-9;
        fc1_weights[103][107] = 16'sd-26;
        fc1_weights[103][108] = 16'sd15;
        fc1_weights[103][109] = 16'sd1;
        fc1_weights[103][110] = 16'sd-26;
        fc1_weights[103][111] = 16'sd57;
        fc1_weights[103][112] = 16'sd-21;
        fc1_weights[103][113] = 16'sd-14;
        fc1_weights[103][114] = 16'sd32;
        fc1_weights[103][115] = 16'sd-9;
        fc1_weights[103][116] = 16'sd37;
        fc1_weights[103][117] = 16'sd34;
        fc1_weights[103][118] = 16'sd48;
        fc1_weights[103][119] = 16'sd30;
        fc1_weights[103][120] = 16'sd-19;
        fc1_weights[103][121] = 16'sd88;
        fc1_weights[103][122] = 16'sd16;
        fc1_weights[103][123] = 16'sd73;
        fc1_weights[103][124] = 16'sd-10;
        fc1_weights[103][125] = 16'sd65;
        fc1_weights[103][126] = 16'sd-43;
        fc1_weights[103][127] = 16'sd21;
        fc1_weights[103][128] = 16'sd41;
        fc1_weights[103][129] = 16'sd-8;
        fc1_weights[103][130] = 16'sd-9;
        fc1_weights[103][131] = 16'sd-27;
        fc1_weights[103][132] = 16'sd-24;
        fc1_weights[103][133] = 16'sd-17;
        fc1_weights[103][134] = 16'sd0;
        fc1_weights[103][135] = 16'sd-7;
        fc1_weights[103][136] = 16'sd12;
        fc1_weights[103][137] = 16'sd36;
        fc1_weights[103][138] = 16'sd45;
        fc1_weights[103][139] = 16'sd-29;
        fc1_weights[103][140] = 16'sd-35;
        fc1_weights[103][141] = 16'sd-70;
        fc1_weights[103][142] = 16'sd35;
        fc1_weights[103][143] = 16'sd-28;
        fc1_weights[103][144] = 16'sd25;
        fc1_weights[103][145] = 16'sd-21;
        fc1_weights[103][146] = 16'sd-9;
        fc1_weights[103][147] = 16'sd-4;
        fc1_weights[103][148] = 16'sd-20;
        fc1_weights[103][149] = 16'sd-2;
        fc1_weights[103][150] = 16'sd44;
        fc1_weights[103][151] = 16'sd15;
        fc1_weights[103][152] = 16'sd-18;
        fc1_weights[103][153] = 16'sd26;
        fc1_weights[103][154] = 16'sd-9;
        fc1_weights[103][155] = 16'sd29;
        fc1_weights[103][156] = 16'sd-9;
        fc1_weights[103][157] = 16'sd-19;
        fc1_weights[103][158] = 16'sd-36;
        fc1_weights[103][159] = 16'sd-3;
        fc1_weights[103][160] = 16'sd17;
        fc1_weights[103][161] = 16'sd-10;
        fc1_weights[103][162] = 16'sd28;
        fc1_weights[103][163] = 16'sd11;
        fc1_weights[103][164] = 16'sd-43;
        fc1_weights[103][165] = 16'sd-34;
        fc1_weights[103][166] = 16'sd31;
        fc1_weights[103][167] = 16'sd-21;
        fc1_weights[103][168] = 16'sd42;
        fc1_weights[103][169] = 16'sd31;
        fc1_weights[103][170] = 16'sd30;
        fc1_weights[103][171] = 16'sd37;
        fc1_weights[103][172] = 16'sd27;
        fc1_weights[103][173] = 16'sd24;
        fc1_weights[103][174] = 16'sd16;
        fc1_weights[103][175] = 16'sd43;
        fc1_weights[103][176] = 16'sd57;
        fc1_weights[103][177] = 16'sd24;
        fc1_weights[103][178] = 16'sd-40;
        fc1_weights[103][179] = 16'sd41;
        fc1_weights[103][180] = 16'sd30;
        fc1_weights[103][181] = 16'sd31;
        fc1_weights[103][182] = 16'sd-20;
        fc1_weights[103][183] = 16'sd-29;
        fc1_weights[103][184] = 16'sd-60;
        fc1_weights[103][185] = 16'sd-10;
        fc1_weights[103][186] = 16'sd-19;
        fc1_weights[103][187] = 16'sd28;
        fc1_weights[103][188] = 16'sd-19;
        fc1_weights[103][189] = 16'sd8;
        fc1_weights[103][190] = 16'sd-63;
        fc1_weights[103][191] = 16'sd5;
        fc1_weights[103][192] = 16'sd-34;
        fc1_weights[103][193] = 16'sd28;
        fc1_weights[103][194] = 16'sd23;
        fc1_weights[103][195] = 16'sd32;
        fc1_weights[103][196] = 16'sd45;
        fc1_weights[103][197] = 16'sd36;
        fc1_weights[103][198] = 16'sd30;
        fc1_weights[103][199] = 16'sd37;
        fc1_weights[103][200] = 16'sd29;
        fc1_weights[103][201] = 16'sd19;
        fc1_weights[103][202] = 16'sd2;
        fc1_weights[103][203] = 16'sd-11;
        fc1_weights[103][204] = 16'sd42;
        fc1_weights[103][205] = 16'sd12;
        fc1_weights[103][206] = 16'sd0;
        fc1_weights[103][207] = 16'sd-46;
        fc1_weights[104][0] = 16'sd26;
        fc1_weights[104][1] = 16'sd8;
        fc1_weights[104][2] = 16'sd15;
        fc1_weights[104][3] = 16'sd-75;
        fc1_weights[104][4] = 16'sd-13;
        fc1_weights[104][5] = 16'sd-22;
        fc1_weights[104][6] = 16'sd-53;
        fc1_weights[104][7] = 16'sd-34;
        fc1_weights[104][8] = 16'sd-82;
        fc1_weights[104][9] = 16'sd36;
        fc1_weights[104][10] = 16'sd10;
        fc1_weights[104][11] = 16'sd-67;
        fc1_weights[104][12] = 16'sd-63;
        fc1_weights[104][13] = 16'sd5;
        fc1_weights[104][14] = 16'sd-5;
        fc1_weights[104][15] = 16'sd65;
        fc1_weights[104][16] = 16'sd-43;
        fc1_weights[104][17] = 16'sd-88;
        fc1_weights[104][18] = 16'sd-22;
        fc1_weights[104][19] = 16'sd-53;
        fc1_weights[104][20] = 16'sd52;
        fc1_weights[104][21] = 16'sd-5;
        fc1_weights[104][22] = 16'sd-31;
        fc1_weights[104][23] = 16'sd-47;
        fc1_weights[104][24] = 16'sd65;
        fc1_weights[104][25] = 16'sd-19;
        fc1_weights[104][26] = 16'sd14;
        fc1_weights[104][27] = 16'sd13;
        fc1_weights[104][28] = 16'sd39;
        fc1_weights[104][29] = 16'sd-26;
        fc1_weights[104][30] = 16'sd-39;
        fc1_weights[104][31] = 16'sd-31;
        fc1_weights[104][32] = 16'sd-51;
        fc1_weights[104][33] = 16'sd-62;
        fc1_weights[104][34] = 16'sd-57;
        fc1_weights[104][35] = 16'sd-25;
        fc1_weights[104][36] = 16'sd49;
        fc1_weights[104][37] = 16'sd-124;
        fc1_weights[104][38] = 16'sd-37;
        fc1_weights[104][39] = 16'sd-31;
        fc1_weights[104][40] = 16'sd42;
        fc1_weights[104][41] = 16'sd19;
        fc1_weights[104][42] = 16'sd-50;
        fc1_weights[104][43] = 16'sd36;
        fc1_weights[104][44] = 16'sd3;
        fc1_weights[104][45] = 16'sd-20;
        fc1_weights[104][46] = 16'sd42;
        fc1_weights[104][47] = 16'sd61;
        fc1_weights[104][48] = 16'sd-28;
        fc1_weights[104][49] = 16'sd20;
        fc1_weights[104][50] = 16'sd43;
        fc1_weights[104][51] = 16'sd-41;
        fc1_weights[104][52] = 16'sd54;
        fc1_weights[104][53] = 16'sd54;
        fc1_weights[104][54] = 16'sd0;
        fc1_weights[104][55] = 16'sd-1;
        fc1_weights[104][56] = 16'sd13;
        fc1_weights[104][57] = 16'sd10;
        fc1_weights[104][58] = 16'sd4;
        fc1_weights[104][59] = 16'sd-2;
        fc1_weights[104][60] = 16'sd30;
        fc1_weights[104][61] = 16'sd19;
        fc1_weights[104][62] = 16'sd-63;
        fc1_weights[104][63] = 16'sd-9;
        fc1_weights[104][64] = 16'sd-12;
        fc1_weights[104][65] = 16'sd-97;
        fc1_weights[104][66] = 16'sd16;
        fc1_weights[104][67] = 16'sd-7;
        fc1_weights[104][68] = 16'sd-4;
        fc1_weights[104][69] = 16'sd-76;
        fc1_weights[104][70] = 16'sd12;
        fc1_weights[104][71] = 16'sd45;
        fc1_weights[104][72] = 16'sd82;
        fc1_weights[104][73] = 16'sd-22;
        fc1_weights[104][74] = 16'sd-59;
        fc1_weights[104][75] = 16'sd-6;
        fc1_weights[104][76] = 16'sd18;
        fc1_weights[104][77] = 16'sd-60;
        fc1_weights[104][78] = 16'sd20;
        fc1_weights[104][79] = 16'sd144;
        fc1_weights[104][80] = 16'sd-5;
        fc1_weights[104][81] = 16'sd3;
        fc1_weights[104][82] = 16'sd10;
        fc1_weights[104][83] = 16'sd10;
        fc1_weights[104][84] = 16'sd-18;
        fc1_weights[104][85] = 16'sd-17;
        fc1_weights[104][86] = 16'sd32;
        fc1_weights[104][87] = 16'sd-16;
        fc1_weights[104][88] = 16'sd19;
        fc1_weights[104][89] = 16'sd-45;
        fc1_weights[104][90] = 16'sd85;
        fc1_weights[104][91] = 16'sd87;
        fc1_weights[104][92] = 16'sd50;
        fc1_weights[104][93] = 16'sd-46;
        fc1_weights[104][94] = 16'sd-50;
        fc1_weights[104][95] = 16'sd-38;
        fc1_weights[104][96] = 16'sd-41;
        fc1_weights[104][97] = 16'sd-56;
        fc1_weights[104][98] = 16'sd-18;
        fc1_weights[104][99] = 16'sd21;
        fc1_weights[104][100] = 16'sd-16;
        fc1_weights[104][101] = 16'sd-86;
        fc1_weights[104][102] = 16'sd-51;
        fc1_weights[104][103] = 16'sd-122;
        fc1_weights[104][104] = 16'sd84;
        fc1_weights[104][105] = 16'sd-10;
        fc1_weights[104][106] = 16'sd12;
        fc1_weights[104][107] = 16'sd42;
        fc1_weights[104][108] = 16'sd-2;
        fc1_weights[104][109] = 16'sd32;
        fc1_weights[104][110] = 16'sd48;
        fc1_weights[104][111] = 16'sd8;
        fc1_weights[104][112] = 16'sd67;
        fc1_weights[104][113] = 16'sd-14;
        fc1_weights[104][114] = 16'sd12;
        fc1_weights[104][115] = 16'sd-33;
        fc1_weights[104][116] = 16'sd13;
        fc1_weights[104][117] = 16'sd27;
        fc1_weights[104][118] = 16'sd11;
        fc1_weights[104][119] = 16'sd15;
        fc1_weights[104][120] = 16'sd-44;
        fc1_weights[104][121] = 16'sd-5;
        fc1_weights[104][122] = 16'sd-29;
        fc1_weights[104][123] = 16'sd-30;
        fc1_weights[104][124] = 16'sd-89;
        fc1_weights[104][125] = 16'sd34;
        fc1_weights[104][126] = 16'sd-105;
        fc1_weights[104][127] = 16'sd-22;
        fc1_weights[104][128] = 16'sd-54;
        fc1_weights[104][129] = 16'sd-130;
        fc1_weights[104][130] = 16'sd14;
        fc1_weights[104][131] = 16'sd27;
        fc1_weights[104][132] = 16'sd36;
        fc1_weights[104][133] = 16'sd5;
        fc1_weights[104][134] = 16'sd-3;
        fc1_weights[104][135] = 16'sd28;
        fc1_weights[104][136] = 16'sd79;
        fc1_weights[104][137] = 16'sd53;
        fc1_weights[104][138] = 16'sd2;
        fc1_weights[104][139] = 16'sd-33;
        fc1_weights[104][140] = 16'sd-35;
        fc1_weights[104][141] = 16'sd-52;
        fc1_weights[104][142] = 16'sd-13;
        fc1_weights[104][143] = 16'sd-3;
        fc1_weights[104][144] = 16'sd-25;
        fc1_weights[104][145] = 16'sd-50;
        fc1_weights[104][146] = 16'sd-15;
        fc1_weights[104][147] = 16'sd70;
        fc1_weights[104][148] = 16'sd51;
        fc1_weights[104][149] = 16'sd-51;
        fc1_weights[104][150] = 16'sd-59;
        fc1_weights[104][151] = 16'sd34;
        fc1_weights[104][152] = 16'sd23;
        fc1_weights[104][153] = 16'sd16;
        fc1_weights[104][154] = 16'sd7;
        fc1_weights[104][155] = 16'sd-3;
        fc1_weights[104][156] = 16'sd3;
        fc1_weights[104][157] = 16'sd71;
        fc1_weights[104][158] = 16'sd27;
        fc1_weights[104][159] = 16'sd21;
        fc1_weights[104][160] = 16'sd-88;
        fc1_weights[104][161] = 16'sd41;
        fc1_weights[104][162] = 16'sd0;
        fc1_weights[104][163] = 16'sd12;
        fc1_weights[104][164] = 16'sd-1;
        fc1_weights[104][165] = 16'sd-75;
        fc1_weights[104][166] = 16'sd-25;
        fc1_weights[104][167] = 16'sd-38;
        fc1_weights[104][168] = 16'sd-91;
        fc1_weights[104][169] = 16'sd25;
        fc1_weights[104][170] = 16'sd47;
        fc1_weights[104][171] = 16'sd44;
        fc1_weights[104][172] = 16'sd7;
        fc1_weights[104][173] = 16'sd26;
        fc1_weights[104][174] = 16'sd0;
        fc1_weights[104][175] = 16'sd40;
        fc1_weights[104][176] = 16'sd-39;
        fc1_weights[104][177] = 16'sd-18;
        fc1_weights[104][178] = 16'sd-2;
        fc1_weights[104][179] = 16'sd1;
        fc1_weights[104][180] = 16'sd10;
        fc1_weights[104][181] = 16'sd49;
        fc1_weights[104][182] = 16'sd12;
        fc1_weights[104][183] = 16'sd63;
        fc1_weights[104][184] = 16'sd2;
        fc1_weights[104][185] = 16'sd66;
        fc1_weights[104][186] = 16'sd-7;
        fc1_weights[104][187] = 16'sd7;
        fc1_weights[104][188] = 16'sd-38;
        fc1_weights[104][189] = 16'sd36;
        fc1_weights[104][190] = 16'sd40;
        fc1_weights[104][191] = 16'sd-35;
        fc1_weights[104][192] = 16'sd-87;
        fc1_weights[104][193] = 16'sd-64;
        fc1_weights[104][194] = 16'sd-41;
        fc1_weights[104][195] = 16'sd-11;
        fc1_weights[104][196] = 16'sd23;
        fc1_weights[104][197] = 16'sd61;
        fc1_weights[104][198] = 16'sd-26;
        fc1_weights[104][199] = 16'sd49;
        fc1_weights[104][200] = 16'sd48;
        fc1_weights[104][201] = 16'sd35;
        fc1_weights[104][202] = 16'sd20;
        fc1_weights[104][203] = 16'sd77;
        fc1_weights[104][204] = 16'sd12;
        fc1_weights[104][205] = 16'sd15;
        fc1_weights[104][206] = 16'sd-63;
        fc1_weights[104][207] = 16'sd-37;
        fc1_weights[105][0] = 16'sd-13;
        fc1_weights[105][1] = 16'sd-10;
        fc1_weights[105][2] = 16'sd24;
        fc1_weights[105][3] = 16'sd-28;
        fc1_weights[105][4] = 16'sd0;
        fc1_weights[105][5] = 16'sd8;
        fc1_weights[105][6] = 16'sd14;
        fc1_weights[105][7] = 16'sd27;
        fc1_weights[105][8] = 16'sd-6;
        fc1_weights[105][9] = 16'sd10;
        fc1_weights[105][10] = 16'sd-12;
        fc1_weights[105][11] = 16'sd-46;
        fc1_weights[105][12] = 16'sd-6;
        fc1_weights[105][13] = 16'sd-24;
        fc1_weights[105][14] = 16'sd-38;
        fc1_weights[105][15] = 16'sd-39;
        fc1_weights[105][16] = 16'sd2;
        fc1_weights[105][17] = 16'sd35;
        fc1_weights[105][18] = 16'sd11;
        fc1_weights[105][19] = 16'sd28;
        fc1_weights[105][20] = 16'sd42;
        fc1_weights[105][21] = 16'sd26;
        fc1_weights[105][22] = 16'sd48;
        fc1_weights[105][23] = 16'sd88;
        fc1_weights[105][24] = 16'sd39;
        fc1_weights[105][25] = 16'sd38;
        fc1_weights[105][26] = 16'sd-11;
        fc1_weights[105][27] = 16'sd-14;
        fc1_weights[105][28] = 16'sd-4;
        fc1_weights[105][29] = 16'sd6;
        fc1_weights[105][30] = 16'sd-16;
        fc1_weights[105][31] = 16'sd23;
        fc1_weights[105][32] = 16'sd8;
        fc1_weights[105][33] = 16'sd31;
        fc1_weights[105][34] = 16'sd14;
        fc1_weights[105][35] = 16'sd-10;
        fc1_weights[105][36] = 16'sd-22;
        fc1_weights[105][37] = 16'sd10;
        fc1_weights[105][38] = 16'sd-20;
        fc1_weights[105][39] = 16'sd-25;
        fc1_weights[105][40] = 16'sd-42;
        fc1_weights[105][41] = 16'sd-28;
        fc1_weights[105][42] = 16'sd-1;
        fc1_weights[105][43] = 16'sd-27;
        fc1_weights[105][44] = 16'sd-26;
        fc1_weights[105][45] = 16'sd-20;
        fc1_weights[105][46] = 16'sd40;
        fc1_weights[105][47] = 16'sd15;
        fc1_weights[105][48] = 16'sd34;
        fc1_weights[105][49] = 16'sd19;
        fc1_weights[105][50] = 16'sd21;
        fc1_weights[105][51] = 16'sd34;
        fc1_weights[105][52] = 16'sd-5;
        fc1_weights[105][53] = 16'sd-24;
        fc1_weights[105][54] = 16'sd-27;
        fc1_weights[105][55] = 16'sd-18;
        fc1_weights[105][56] = 16'sd-27;
        fc1_weights[105][57] = 16'sd-27;
        fc1_weights[105][58] = 16'sd-34;
        fc1_weights[105][59] = 16'sd-42;
        fc1_weights[105][60] = 16'sd-49;
        fc1_weights[105][61] = 16'sd-43;
        fc1_weights[105][62] = 16'sd-10;
        fc1_weights[105][63] = 16'sd-4;
        fc1_weights[105][64] = 16'sd-27;
        fc1_weights[105][65] = 16'sd-36;
        fc1_weights[105][66] = 16'sd-28;
        fc1_weights[105][67] = 16'sd-17;
        fc1_weights[105][68] = 16'sd0;
        fc1_weights[105][69] = 16'sd33;
        fc1_weights[105][70] = 16'sd15;
        fc1_weights[105][71] = 16'sd29;
        fc1_weights[105][72] = 16'sd23;
        fc1_weights[105][73] = 16'sd40;
        fc1_weights[105][74] = 16'sd9;
        fc1_weights[105][75] = 16'sd34;
        fc1_weights[105][76] = 16'sd1;
        fc1_weights[105][77] = 16'sd1;
        fc1_weights[105][78] = 16'sd-25;
        fc1_weights[105][79] = 16'sd-8;
        fc1_weights[105][80] = 16'sd-6;
        fc1_weights[105][81] = 16'sd17;
        fc1_weights[105][82] = 16'sd-18;
        fc1_weights[105][83] = 16'sd-18;
        fc1_weights[105][84] = 16'sd6;
        fc1_weights[105][85] = 16'sd8;
        fc1_weights[105][86] = 16'sd6;
        fc1_weights[105][87] = 16'sd8;
        fc1_weights[105][88] = 16'sd-16;
        fc1_weights[105][89] = 16'sd2;
        fc1_weights[105][90] = 16'sd-41;
        fc1_weights[105][91] = 16'sd-33;
        fc1_weights[105][92] = 16'sd-27;
        fc1_weights[105][93] = 16'sd25;
        fc1_weights[105][94] = 16'sd25;
        fc1_weights[105][95] = 16'sd23;
        fc1_weights[105][96] = 16'sd21;
        fc1_weights[105][97] = 16'sd-13;
        fc1_weights[105][98] = 16'sd10;
        fc1_weights[105][99] = 16'sd24;
        fc1_weights[105][100] = 16'sd38;
        fc1_weights[105][101] = 16'sd29;
        fc1_weights[105][102] = 16'sd11;
        fc1_weights[105][103] = 16'sd20;
        fc1_weights[105][104] = 16'sd-26;
        fc1_weights[105][105] = 16'sd-22;
        fc1_weights[105][106] = 16'sd-15;
        fc1_weights[105][107] = 16'sd-16;
        fc1_weights[105][108] = 16'sd-18;
        fc1_weights[105][109] = 16'sd-13;
        fc1_weights[105][110] = 16'sd8;
        fc1_weights[105][111] = 16'sd7;
        fc1_weights[105][112] = 16'sd-40;
        fc1_weights[105][113] = 16'sd-33;
        fc1_weights[105][114] = 16'sd-21;
        fc1_weights[105][115] = 16'sd6;
        fc1_weights[105][116] = 16'sd-19;
        fc1_weights[105][117] = 16'sd-7;
        fc1_weights[105][118] = 16'sd-20;
        fc1_weights[105][119] = 16'sd0;
        fc1_weights[105][120] = 16'sd5;
        fc1_weights[105][121] = 16'sd19;
        fc1_weights[105][122] = 16'sd39;
        fc1_weights[105][123] = 16'sd-8;
        fc1_weights[105][124] = 16'sd57;
        fc1_weights[105][125] = 16'sd23;
        fc1_weights[105][126] = 16'sd31;
        fc1_weights[105][127] = 16'sd26;
        fc1_weights[105][128] = 16'sd49;
        fc1_weights[105][129] = 16'sd77;
        fc1_weights[105][130] = 16'sd-8;
        fc1_weights[105][131] = 16'sd5;
        fc1_weights[105][132] = 16'sd3;
        fc1_weights[105][133] = 16'sd-2;
        fc1_weights[105][134] = 16'sd-27;
        fc1_weights[105][135] = 16'sd-20;
        fc1_weights[105][136] = 16'sd3;
        fc1_weights[105][137] = 16'sd-4;
        fc1_weights[105][138] = 16'sd-37;
        fc1_weights[105][139] = 16'sd2;
        fc1_weights[105][140] = 16'sd13;
        fc1_weights[105][141] = 16'sd30;
        fc1_weights[105][142] = 16'sd8;
        fc1_weights[105][143] = 16'sd8;
        fc1_weights[105][144] = 16'sd-21;
        fc1_weights[105][145] = 16'sd0;
        fc1_weights[105][146] = 16'sd-10;
        fc1_weights[105][147] = 16'sd-24;
        fc1_weights[105][148] = 16'sd4;
        fc1_weights[105][149] = 16'sd3;
        fc1_weights[105][150] = 16'sd28;
        fc1_weights[105][151] = 16'sd8;
        fc1_weights[105][152] = 16'sd21;
        fc1_weights[105][153] = 16'sd27;
        fc1_weights[105][154] = 16'sd19;
        fc1_weights[105][155] = 16'sd6;
        fc1_weights[105][156] = 16'sd14;
        fc1_weights[105][157] = 16'sd7;
        fc1_weights[105][158] = 16'sd12;
        fc1_weights[105][159] = 16'sd9;
        fc1_weights[105][160] = 16'sd27;
        fc1_weights[105][161] = 16'sd-4;
        fc1_weights[105][162] = 16'sd-15;
        fc1_weights[105][163] = 16'sd29;
        fc1_weights[105][164] = 16'sd39;
        fc1_weights[105][165] = 16'sd7;
        fc1_weights[105][166] = 16'sd14;
        fc1_weights[105][167] = 16'sd-13;
        fc1_weights[105][168] = 16'sd7;
        fc1_weights[105][169] = 16'sd4;
        fc1_weights[105][170] = 16'sd-14;
        fc1_weights[105][171] = 16'sd-21;
        fc1_weights[105][172] = 16'sd-13;
        fc1_weights[105][173] = 16'sd-20;
        fc1_weights[105][174] = 16'sd10;
        fc1_weights[105][175] = 16'sd15;
        fc1_weights[105][176] = 16'sd13;
        fc1_weights[105][177] = 16'sd3;
        fc1_weights[105][178] = 16'sd22;
        fc1_weights[105][179] = 16'sd14;
        fc1_weights[105][180] = 16'sd20;
        fc1_weights[105][181] = 16'sd10;
        fc1_weights[105][182] = 16'sd8;
        fc1_weights[105][183] = 16'sd-8;
        fc1_weights[105][184] = 16'sd-15;
        fc1_weights[105][185] = 16'sd-29;
        fc1_weights[105][186] = 16'sd2;
        fc1_weights[105][187] = 16'sd0;
        fc1_weights[105][188] = 16'sd13;
        fc1_weights[105][189] = 16'sd11;
        fc1_weights[105][190] = 16'sd-8;
        fc1_weights[105][191] = 16'sd-13;
        fc1_weights[105][192] = 16'sd9;
        fc1_weights[105][193] = 16'sd-5;
        fc1_weights[105][194] = 16'sd-9;
        fc1_weights[105][195] = 16'sd-4;
        fc1_weights[105][196] = 16'sd-11;
        fc1_weights[105][197] = 16'sd-22;
        fc1_weights[105][198] = 16'sd-3;
        fc1_weights[105][199] = 16'sd-16;
        fc1_weights[105][200] = 16'sd2;
        fc1_weights[105][201] = 16'sd-1;
        fc1_weights[105][202] = 16'sd23;
        fc1_weights[105][203] = 16'sd-12;
        fc1_weights[105][204] = 16'sd32;
        fc1_weights[105][205] = 16'sd31;
        fc1_weights[105][206] = 16'sd38;
        fc1_weights[105][207] = 16'sd25;
        fc1_weights[106][0] = 16'sd18;
        fc1_weights[106][1] = 16'sd40;
        fc1_weights[106][2] = 16'sd-13;
        fc1_weights[106][3] = 16'sd8;
        fc1_weights[106][4] = 16'sd-4;
        fc1_weights[106][5] = 16'sd21;
        fc1_weights[106][6] = 16'sd29;
        fc1_weights[106][7] = 16'sd23;
        fc1_weights[106][8] = 16'sd-13;
        fc1_weights[106][9] = 16'sd-13;
        fc1_weights[106][10] = 16'sd28;
        fc1_weights[106][11] = 16'sd35;
        fc1_weights[106][12] = 16'sd6;
        fc1_weights[106][13] = 16'sd-3;
        fc1_weights[106][14] = 16'sd15;
        fc1_weights[106][15] = 16'sd17;
        fc1_weights[106][16] = 16'sd45;
        fc1_weights[106][17] = 16'sd26;
        fc1_weights[106][18] = 16'sd4;
        fc1_weights[106][19] = 16'sd0;
        fc1_weights[106][20] = 16'sd20;
        fc1_weights[106][21] = 16'sd22;
        fc1_weights[106][22] = 16'sd1;
        fc1_weights[106][23] = 16'sd26;
        fc1_weights[106][24] = 16'sd-31;
        fc1_weights[106][25] = 16'sd-1;
        fc1_weights[106][26] = 16'sd4;
        fc1_weights[106][27] = 16'sd5;
        fc1_weights[106][28] = 16'sd18;
        fc1_weights[106][29] = 16'sd12;
        fc1_weights[106][30] = 16'sd32;
        fc1_weights[106][31] = 16'sd36;
        fc1_weights[106][32] = 16'sd19;
        fc1_weights[106][33] = 16'sd0;
        fc1_weights[106][34] = 16'sd5;
        fc1_weights[106][35] = 16'sd-2;
        fc1_weights[106][36] = 16'sd7;
        fc1_weights[106][37] = 16'sd27;
        fc1_weights[106][38] = 16'sd26;
        fc1_weights[106][39] = 16'sd-5;
        fc1_weights[106][40] = 16'sd36;
        fc1_weights[106][41] = 16'sd9;
        fc1_weights[106][42] = 16'sd19;
        fc1_weights[106][43] = 16'sd-1;
        fc1_weights[106][44] = 16'sd-2;
        fc1_weights[106][45] = 16'sd1;
        fc1_weights[106][46] = 16'sd-26;
        fc1_weights[106][47] = 16'sd-10;
        fc1_weights[106][48] = 16'sd9;
        fc1_weights[106][49] = 16'sd-14;
        fc1_weights[106][50] = 16'sd-13;
        fc1_weights[106][51] = 16'sd-13;
        fc1_weights[106][52] = 16'sd48;
        fc1_weights[106][53] = 16'sd26;
        fc1_weights[106][54] = 16'sd19;
        fc1_weights[106][55] = 16'sd31;
        fc1_weights[106][56] = 16'sd12;
        fc1_weights[106][57] = 16'sd6;
        fc1_weights[106][58] = 16'sd12;
        fc1_weights[106][59] = 16'sd2;
        fc1_weights[106][60] = 16'sd-10;
        fc1_weights[106][61] = 16'sd-7;
        fc1_weights[106][62] = 16'sd11;
        fc1_weights[106][63] = 16'sd4;
        fc1_weights[106][64] = 16'sd4;
        fc1_weights[106][65] = 16'sd1;
        fc1_weights[106][66] = 16'sd17;
        fc1_weights[106][67] = 16'sd15;
        fc1_weights[106][68] = 16'sd-1;
        fc1_weights[106][69] = 16'sd30;
        fc1_weights[106][70] = 16'sd39;
        fc1_weights[106][71] = 16'sd0;
        fc1_weights[106][72] = 16'sd-14;
        fc1_weights[106][73] = 16'sd1;
        fc1_weights[106][74] = 16'sd-3;
        fc1_weights[106][75] = 16'sd13;
        fc1_weights[106][76] = 16'sd12;
        fc1_weights[106][77] = 16'sd4;
        fc1_weights[106][78] = 16'sd25;
        fc1_weights[106][79] = 16'sd-14;
        fc1_weights[106][80] = 16'sd-2;
        fc1_weights[106][81] = 16'sd0;
        fc1_weights[106][82] = 16'sd1;
        fc1_weights[106][83] = 16'sd32;
        fc1_weights[106][84] = 16'sd27;
        fc1_weights[106][85] = 16'sd16;
        fc1_weights[106][86] = 16'sd-7;
        fc1_weights[106][87] = 16'sd-12;
        fc1_weights[106][88] = 16'sd-18;
        fc1_weights[106][89] = 16'sd-14;
        fc1_weights[106][90] = 16'sd-21;
        fc1_weights[106][91] = 16'sd-14;
        fc1_weights[106][92] = 16'sd2;
        fc1_weights[106][93] = 16'sd15;
        fc1_weights[106][94] = 16'sd8;
        fc1_weights[106][95] = 16'sd0;
        fc1_weights[106][96] = 16'sd24;
        fc1_weights[106][97] = 16'sd4;
        fc1_weights[106][98] = 16'sd-2;
        fc1_weights[106][99] = 16'sd2;
        fc1_weights[106][100] = 16'sd-11;
        fc1_weights[106][101] = 16'sd13;
        fc1_weights[106][102] = 16'sd3;
        fc1_weights[106][103] = 16'sd4;
        fc1_weights[106][104] = 16'sd-4;
        fc1_weights[106][105] = 16'sd-4;
        fc1_weights[106][106] = 16'sd-2;
        fc1_weights[106][107] = 16'sd-16;
        fc1_weights[106][108] = 16'sd-2;
        fc1_weights[106][109] = 16'sd6;
        fc1_weights[106][110] = 16'sd-34;
        fc1_weights[106][111] = 16'sd0;
        fc1_weights[106][112] = 16'sd1;
        fc1_weights[106][113] = 16'sd-18;
        fc1_weights[106][114] = 16'sd-21;
        fc1_weights[106][115] = 16'sd-13;
        fc1_weights[106][116] = 16'sd-38;
        fc1_weights[106][117] = 16'sd-11;
        fc1_weights[106][118] = 16'sd-6;
        fc1_weights[106][119] = 16'sd-4;
        fc1_weights[106][120] = 16'sd15;
        fc1_weights[106][121] = 16'sd16;
        fc1_weights[106][122] = 16'sd6;
        fc1_weights[106][123] = 16'sd-6;
        fc1_weights[106][124] = 16'sd16;
        fc1_weights[106][125] = 16'sd7;
        fc1_weights[106][126] = 16'sd2;
        fc1_weights[106][127] = 16'sd29;
        fc1_weights[106][128] = 16'sd-1;
        fc1_weights[106][129] = 16'sd-5;
        fc1_weights[106][130] = 16'sd-16;
        fc1_weights[106][131] = 16'sd-15;
        fc1_weights[106][132] = 16'sd-26;
        fc1_weights[106][133] = 16'sd-12;
        fc1_weights[106][134] = 16'sd8;
        fc1_weights[106][135] = 16'sd16;
        fc1_weights[106][136] = 16'sd-8;
        fc1_weights[106][137] = 16'sd-13;
        fc1_weights[106][138] = 16'sd24;
        fc1_weights[106][139] = 16'sd33;
        fc1_weights[106][140] = 16'sd-3;
        fc1_weights[106][141] = 16'sd8;
        fc1_weights[106][142] = 16'sd1;
        fc1_weights[106][143] = 16'sd-35;
        fc1_weights[106][144] = 16'sd15;
        fc1_weights[106][145] = 16'sd2;
        fc1_weights[106][146] = 16'sd-16;
        fc1_weights[106][147] = 16'sd-15;
        fc1_weights[106][148] = 16'sd5;
        fc1_weights[106][149] = 16'sd5;
        fc1_weights[106][150] = 16'sd32;
        fc1_weights[106][151] = 16'sd-14;
        fc1_weights[106][152] = 16'sd-5;
        fc1_weights[106][153] = 16'sd-34;
        fc1_weights[106][154] = 16'sd-16;
        fc1_weights[106][155] = 16'sd-19;
        fc1_weights[106][156] = 16'sd-20;
        fc1_weights[106][157] = 16'sd-6;
        fc1_weights[106][158] = 16'sd-21;
        fc1_weights[106][159] = 16'sd-23;
        fc1_weights[106][160] = 16'sd22;
        fc1_weights[106][161] = 16'sd5;
        fc1_weights[106][162] = 16'sd12;
        fc1_weights[106][163] = 16'sd7;
        fc1_weights[106][164] = 16'sd17;
        fc1_weights[106][165] = 16'sd26;
        fc1_weights[106][166] = 16'sd8;
        fc1_weights[106][167] = 16'sd-1;
        fc1_weights[106][168] = 16'sd3;
        fc1_weights[106][169] = 16'sd-10;
        fc1_weights[106][170] = 16'sd-36;
        fc1_weights[106][171] = 16'sd-23;
        fc1_weights[106][172] = 16'sd-18;
        fc1_weights[106][173] = 16'sd-4;
        fc1_weights[106][174] = 16'sd-14;
        fc1_weights[106][175] = 16'sd-28;
        fc1_weights[106][176] = 16'sd-18;
        fc1_weights[106][177] = 16'sd-30;
        fc1_weights[106][178] = 16'sd-14;
        fc1_weights[106][179] = 16'sd-22;
        fc1_weights[106][180] = 16'sd-16;
        fc1_weights[106][181] = 16'sd-13;
        fc1_weights[106][182] = 16'sd1;
        fc1_weights[106][183] = 16'sd-4;
        fc1_weights[106][184] = 16'sd-14;
        fc1_weights[106][185] = 16'sd-27;
        fc1_weights[106][186] = 16'sd30;
        fc1_weights[106][187] = 16'sd23;
        fc1_weights[106][188] = 16'sd7;
        fc1_weights[106][189] = 16'sd10;
        fc1_weights[106][190] = 16'sd21;
        fc1_weights[106][191] = 16'sd17;
        fc1_weights[106][192] = 16'sd32;
        fc1_weights[106][193] = 16'sd17;
        fc1_weights[106][194] = 16'sd0;
        fc1_weights[106][195] = 16'sd5;
        fc1_weights[106][196] = 16'sd-23;
        fc1_weights[106][197] = 16'sd-8;
        fc1_weights[106][198] = 16'sd-16;
        fc1_weights[106][199] = 16'sd-16;
        fc1_weights[106][200] = 16'sd-30;
        fc1_weights[106][201] = 16'sd-29;
        fc1_weights[106][202] = 16'sd-32;
        fc1_weights[106][203] = 16'sd1;
        fc1_weights[106][204] = 16'sd14;
        fc1_weights[106][205] = 16'sd-20;
        fc1_weights[106][206] = 16'sd-18;
        fc1_weights[106][207] = 16'sd-11;
        fc1_weights[107][0] = 16'sd25;
        fc1_weights[107][1] = 16'sd2;
        fc1_weights[107][2] = 16'sd-44;
        fc1_weights[107][3] = 16'sd-68;
        fc1_weights[107][4] = 16'sd-65;
        fc1_weights[107][5] = 16'sd-32;
        fc1_weights[107][6] = 16'sd-63;
        fc1_weights[107][7] = 16'sd-35;
        fc1_weights[107][8] = 16'sd-11;
        fc1_weights[107][9] = 16'sd-18;
        fc1_weights[107][10] = 16'sd36;
        fc1_weights[107][11] = 16'sd-27;
        fc1_weights[107][12] = 16'sd-43;
        fc1_weights[107][13] = 16'sd-32;
        fc1_weights[107][14] = 16'sd0;
        fc1_weights[107][15] = 16'sd39;
        fc1_weights[107][16] = 16'sd18;
        fc1_weights[107][17] = 16'sd10;
        fc1_weights[107][18] = 16'sd33;
        fc1_weights[107][19] = 16'sd-9;
        fc1_weights[107][20] = 16'sd20;
        fc1_weights[107][21] = 16'sd39;
        fc1_weights[107][22] = 16'sd12;
        fc1_weights[107][23] = 16'sd-19;
        fc1_weights[107][24] = 16'sd44;
        fc1_weights[107][25] = 16'sd44;
        fc1_weights[107][26] = 16'sd32;
        fc1_weights[107][27] = 16'sd-46;
        fc1_weights[107][28] = 16'sd-49;
        fc1_weights[107][29] = 16'sd-21;
        fc1_weights[107][30] = 16'sd5;
        fc1_weights[107][31] = 16'sd16;
        fc1_weights[107][32] = 16'sd-24;
        fc1_weights[107][33] = 16'sd-87;
        fc1_weights[107][34] = 16'sd-22;
        fc1_weights[107][35] = 16'sd1;
        fc1_weights[107][36] = 16'sd25;
        fc1_weights[107][37] = 16'sd37;
        fc1_weights[107][38] = 16'sd-29;
        fc1_weights[107][39] = 16'sd-47;
        fc1_weights[107][40] = 16'sd31;
        fc1_weights[107][41] = 16'sd27;
        fc1_weights[107][42] = 16'sd16;
        fc1_weights[107][43] = 16'sd16;
        fc1_weights[107][44] = 16'sd-6;
        fc1_weights[107][45] = 16'sd-29;
        fc1_weights[107][46] = 16'sd-40;
        fc1_weights[107][47] = 16'sd16;
        fc1_weights[107][48] = 16'sd-1;
        fc1_weights[107][49] = 16'sd-1;
        fc1_weights[107][50] = 16'sd68;
        fc1_weights[107][51] = 16'sd-3;
        fc1_weights[107][52] = 16'sd1;
        fc1_weights[107][53] = 16'sd70;
        fc1_weights[107][54] = 16'sd-25;
        fc1_weights[107][55] = 16'sd45;
        fc1_weights[107][56] = 16'sd9;
        fc1_weights[107][57] = 16'sd56;
        fc1_weights[107][58] = 16'sd65;
        fc1_weights[107][59] = 16'sd11;
        fc1_weights[107][60] = 16'sd-30;
        fc1_weights[107][61] = 16'sd6;
        fc1_weights[107][62] = 16'sd-24;
        fc1_weights[107][63] = 16'sd20;
        fc1_weights[107][64] = 16'sd-21;
        fc1_weights[107][65] = 16'sd-25;
        fc1_weights[107][66] = 16'sd-6;
        fc1_weights[107][67] = 16'sd18;
        fc1_weights[107][68] = 16'sd-13;
        fc1_weights[107][69] = 16'sd-12;
        fc1_weights[107][70] = 16'sd13;
        fc1_weights[107][71] = 16'sd-44;
        fc1_weights[107][72] = 16'sd-24;
        fc1_weights[107][73] = 16'sd13;
        fc1_weights[107][74] = 16'sd-52;
        fc1_weights[107][75] = 16'sd-32;
        fc1_weights[107][76] = 16'sd-22;
        fc1_weights[107][77] = 16'sd-45;
        fc1_weights[107][78] = 16'sd-25;
        fc1_weights[107][79] = 16'sd24;
        fc1_weights[107][80] = 16'sd49;
        fc1_weights[107][81] = 16'sd22;
        fc1_weights[107][82] = 16'sd28;
        fc1_weights[107][83] = 16'sd41;
        fc1_weights[107][84] = 16'sd11;
        fc1_weights[107][85] = 16'sd-50;
        fc1_weights[107][86] = 16'sd-8;
        fc1_weights[107][87] = 16'sd-35;
        fc1_weights[107][88] = 16'sd2;
        fc1_weights[107][89] = 16'sd-4;
        fc1_weights[107][90] = 16'sd-54;
        fc1_weights[107][91] = 16'sd-60;
        fc1_weights[107][92] = 16'sd-13;
        fc1_weights[107][93] = 16'sd49;
        fc1_weights[107][94] = 16'sd-24;
        fc1_weights[107][95] = 16'sd-37;
        fc1_weights[107][96] = 16'sd-13;
        fc1_weights[107][97] = 16'sd-16;
        fc1_weights[107][98] = 16'sd-7;
        fc1_weights[107][99] = 16'sd19;
        fc1_weights[107][100] = 16'sd-37;
        fc1_weights[107][101] = 16'sd-75;
        fc1_weights[107][102] = 16'sd-53;
        fc1_weights[107][103] = 16'sd-39;
        fc1_weights[107][104] = 16'sd34;
        fc1_weights[107][105] = 16'sd-1;
        fc1_weights[107][106] = 16'sd78;
        fc1_weights[107][107] = 16'sd10;
        fc1_weights[107][108] = 16'sd72;
        fc1_weights[107][109] = 16'sd16;
        fc1_weights[107][110] = 16'sd83;
        fc1_weights[107][111] = 16'sd-51;
        fc1_weights[107][112] = 16'sd29;
        fc1_weights[107][113] = 16'sd57;
        fc1_weights[107][114] = 16'sd-7;
        fc1_weights[107][115] = 16'sd40;
        fc1_weights[107][116] = 16'sd-57;
        fc1_weights[107][117] = 16'sd18;
        fc1_weights[107][118] = 16'sd-3;
        fc1_weights[107][119] = 16'sd-3;
        fc1_weights[107][120] = 16'sd-33;
        fc1_weights[107][121] = 16'sd-15;
        fc1_weights[107][122] = 16'sd-1;
        fc1_weights[107][123] = 16'sd-23;
        fc1_weights[107][124] = 16'sd-67;
        fc1_weights[107][125] = 16'sd-64;
        fc1_weights[107][126] = 16'sd-46;
        fc1_weights[107][127] = 16'sd11;
        fc1_weights[107][128] = 16'sd-59;
        fc1_weights[107][129] = 16'sd-85;
        fc1_weights[107][130] = 16'sd12;
        fc1_weights[107][131] = 16'sd-35;
        fc1_weights[107][132] = 16'sd7;
        fc1_weights[107][133] = 16'sd-6;
        fc1_weights[107][134] = 16'sd-20;
        fc1_weights[107][135] = 16'sd-8;
        fc1_weights[107][136] = 16'sd-7;
        fc1_weights[107][137] = 16'sd-6;
        fc1_weights[107][138] = 16'sd55;
        fc1_weights[107][139] = 16'sd35;
        fc1_weights[107][140] = 16'sd25;
        fc1_weights[107][141] = 16'sd57;
        fc1_weights[107][142] = 16'sd-37;
        fc1_weights[107][143] = 16'sd4;
        fc1_weights[107][144] = 16'sd53;
        fc1_weights[107][145] = 16'sd27;
        fc1_weights[107][146] = 16'sd-17;
        fc1_weights[107][147] = 16'sd34;
        fc1_weights[107][148] = 16'sd0;
        fc1_weights[107][149] = 16'sd-32;
        fc1_weights[107][150] = 16'sd-25;
        fc1_weights[107][151] = 16'sd-10;
        fc1_weights[107][152] = 16'sd-24;
        fc1_weights[107][153] = 16'sd14;
        fc1_weights[107][154] = 16'sd-21;
        fc1_weights[107][155] = 16'sd37;
        fc1_weights[107][156] = 16'sd-22;
        fc1_weights[107][157] = 16'sd17;
        fc1_weights[107][158] = 16'sd-34;
        fc1_weights[107][159] = 16'sd-3;
        fc1_weights[107][160] = 16'sd-5;
        fc1_weights[107][161] = 16'sd-15;
        fc1_weights[107][162] = 16'sd19;
        fc1_weights[107][163] = 16'sd12;
        fc1_weights[107][164] = 16'sd11;
        fc1_weights[107][165] = 16'sd25;
        fc1_weights[107][166] = 16'sd-4;
        fc1_weights[107][167] = 16'sd12;
        fc1_weights[107][168] = 16'sd7;
        fc1_weights[107][169] = 16'sd11;
        fc1_weights[107][170] = 16'sd49;
        fc1_weights[107][171] = 16'sd22;
        fc1_weights[107][172] = 16'sd86;
        fc1_weights[107][173] = 16'sd37;
        fc1_weights[107][174] = 16'sd14;
        fc1_weights[107][175] = 16'sd-26;
        fc1_weights[107][176] = 16'sd-12;
        fc1_weights[107][177] = 16'sd21;
        fc1_weights[107][178] = 16'sd0;
        fc1_weights[107][179] = 16'sd19;
        fc1_weights[107][180] = 16'sd32;
        fc1_weights[107][181] = 16'sd1;
        fc1_weights[107][182] = 16'sd-9;
        fc1_weights[107][183] = 16'sd-28;
        fc1_weights[107][184] = 16'sd-24;
        fc1_weights[107][185] = 16'sd34;
        fc1_weights[107][186] = 16'sd27;
        fc1_weights[107][187] = 16'sd8;
        fc1_weights[107][188] = 16'sd13;
        fc1_weights[107][189] = 16'sd11;
        fc1_weights[107][190] = 16'sd38;
        fc1_weights[107][191] = 16'sd2;
        fc1_weights[107][192] = 16'sd8;
        fc1_weights[107][193] = 16'sd2;
        fc1_weights[107][194] = 16'sd-28;
        fc1_weights[107][195] = 16'sd5;
        fc1_weights[107][196] = 16'sd4;
        fc1_weights[107][197] = 16'sd16;
        fc1_weights[107][198] = 16'sd-16;
        fc1_weights[107][199] = 16'sd83;
        fc1_weights[107][200] = 16'sd63;
        fc1_weights[107][201] = 16'sd29;
        fc1_weights[107][202] = 16'sd24;
        fc1_weights[107][203] = 16'sd81;
        fc1_weights[107][204] = 16'sd43;
        fc1_weights[107][205] = 16'sd22;
        fc1_weights[107][206] = 16'sd20;
        fc1_weights[107][207] = 16'sd-14;
        fc1_weights[108][0] = 16'sd47;
        fc1_weights[108][1] = 16'sd50;
        fc1_weights[108][2] = 16'sd1;
        fc1_weights[108][3] = 16'sd44;
        fc1_weights[108][4] = 16'sd34;
        fc1_weights[108][5] = 16'sd12;
        fc1_weights[108][6] = 16'sd0;
        fc1_weights[108][7] = 16'sd88;
        fc1_weights[108][8] = 16'sd-5;
        fc1_weights[108][9] = 16'sd-16;
        fc1_weights[108][10] = 16'sd-6;
        fc1_weights[108][11] = 16'sd14;
        fc1_weights[108][12] = 16'sd13;
        fc1_weights[108][13] = 16'sd-77;
        fc1_weights[108][14] = 16'sd-4;
        fc1_weights[108][15] = 16'sd-46;
        fc1_weights[108][16] = 16'sd2;
        fc1_weights[108][17] = 16'sd8;
        fc1_weights[108][18] = 16'sd18;
        fc1_weights[108][19] = 16'sd34;
        fc1_weights[108][20] = 16'sd62;
        fc1_weights[108][21] = 16'sd35;
        fc1_weights[108][22] = 16'sd2;
        fc1_weights[108][23] = 16'sd25;
        fc1_weights[108][24] = 16'sd10;
        fc1_weights[108][25] = 16'sd-29;
        fc1_weights[108][26] = 16'sd-21;
        fc1_weights[108][27] = 16'sd5;
        fc1_weights[108][28] = 16'sd0;
        fc1_weights[108][29] = 16'sd6;
        fc1_weights[108][30] = 16'sd-10;
        fc1_weights[108][31] = 16'sd-13;
        fc1_weights[108][32] = 16'sd-48;
        fc1_weights[108][33] = 16'sd108;
        fc1_weights[108][34] = 16'sd31;
        fc1_weights[108][35] = 16'sd10;
        fc1_weights[108][36] = 16'sd-3;
        fc1_weights[108][37] = 16'sd54;
        fc1_weights[108][38] = 16'sd46;
        fc1_weights[108][39] = 16'sd-21;
        fc1_weights[108][40] = 16'sd-31;
        fc1_weights[108][41] = 16'sd-29;
        fc1_weights[108][42] = 16'sd16;
        fc1_weights[108][43] = 16'sd-1;
        fc1_weights[108][44] = 16'sd6;
        fc1_weights[108][45] = 16'sd-17;
        fc1_weights[108][46] = 16'sd-21;
        fc1_weights[108][47] = 16'sd31;
        fc1_weights[108][48] = 16'sd4;
        fc1_weights[108][49] = 16'sd-67;
        fc1_weights[108][50] = 16'sd-11;
        fc1_weights[108][51] = 16'sd-16;
        fc1_weights[108][52] = 16'sd-12;
        fc1_weights[108][53] = 16'sd-12;
        fc1_weights[108][54] = 16'sd6;
        fc1_weights[108][55] = 16'sd-10;
        fc1_weights[108][56] = 16'sd-43;
        fc1_weights[108][57] = 16'sd-18;
        fc1_weights[108][58] = 16'sd-6;
        fc1_weights[108][59] = 16'sd20;
        fc1_weights[108][60] = 16'sd-17;
        fc1_weights[108][61] = 16'sd30;
        fc1_weights[108][62] = 16'sd39;
        fc1_weights[108][63] = 16'sd-1;
        fc1_weights[108][64] = 16'sd15;
        fc1_weights[108][65] = 16'sd41;
        fc1_weights[108][66] = 16'sd1;
        fc1_weights[108][67] = 16'sd-36;
        fc1_weights[108][68] = 16'sd-32;
        fc1_weights[108][69] = 16'sd1;
        fc1_weights[108][70] = 16'sd7;
        fc1_weights[108][71] = 16'sd-27;
        fc1_weights[108][72] = 16'sd25;
        fc1_weights[108][73] = 16'sd-10;
        fc1_weights[108][74] = 16'sd-10;
        fc1_weights[108][75] = 16'sd2;
        fc1_weights[108][76] = 16'sd-38;
        fc1_weights[108][77] = 16'sd-15;
        fc1_weights[108][78] = 16'sd-21;
        fc1_weights[108][79] = 16'sd-31;
        fc1_weights[108][80] = 16'sd-3;
        fc1_weights[108][81] = 16'sd-74;
        fc1_weights[108][82] = 16'sd-7;
        fc1_weights[108][83] = 16'sd16;
        fc1_weights[108][84] = 16'sd59;
        fc1_weights[108][85] = 16'sd15;
        fc1_weights[108][86] = 16'sd-24;
        fc1_weights[108][87] = 16'sd-33;
        fc1_weights[108][88] = 16'sd-21;
        fc1_weights[108][89] = 16'sd-48;
        fc1_weights[108][90] = 16'sd5;
        fc1_weights[108][91] = 16'sd-45;
        fc1_weights[108][92] = 16'sd-67;
        fc1_weights[108][93] = 16'sd-30;
        fc1_weights[108][94] = 16'sd3;
        fc1_weights[108][95] = 16'sd-12;
        fc1_weights[108][96] = 16'sd5;
        fc1_weights[108][97] = 16'sd-1;
        fc1_weights[108][98] = 16'sd0;
        fc1_weights[108][99] = 16'sd-24;
        fc1_weights[108][100] = 16'sd19;
        fc1_weights[108][101] = 16'sd49;
        fc1_weights[108][102] = 16'sd28;
        fc1_weights[108][103] = 16'sd17;
        fc1_weights[108][104] = 16'sd-8;
        fc1_weights[108][105] = 16'sd33;
        fc1_weights[108][106] = 16'sd-38;
        fc1_weights[108][107] = 16'sd-47;
        fc1_weights[108][108] = 16'sd-26;
        fc1_weights[108][109] = 16'sd-4;
        fc1_weights[108][110] = 16'sd1;
        fc1_weights[108][111] = 16'sd3;
        fc1_weights[108][112] = 16'sd-35;
        fc1_weights[108][113] = 16'sd3;
        fc1_weights[108][114] = 16'sd-10;
        fc1_weights[108][115] = 16'sd-18;
        fc1_weights[108][116] = 16'sd35;
        fc1_weights[108][117] = 16'sd-40;
        fc1_weights[108][118] = 16'sd-68;
        fc1_weights[108][119] = 16'sd-113;
        fc1_weights[108][120] = 16'sd-60;
        fc1_weights[108][121] = 16'sd-55;
        fc1_weights[108][122] = 16'sd0;
        fc1_weights[108][123] = 16'sd-82;
        fc1_weights[108][124] = 16'sd-12;
        fc1_weights[108][125] = 16'sd-46;
        fc1_weights[108][126] = 16'sd-21;
        fc1_weights[108][127] = 16'sd-55;
        fc1_weights[108][128] = 16'sd-37;
        fc1_weights[108][129] = 16'sd-8;
        fc1_weights[108][130] = 16'sd50;
        fc1_weights[108][131] = 16'sd-21;
        fc1_weights[108][132] = 16'sd-24;
        fc1_weights[108][133] = 16'sd-1;
        fc1_weights[108][134] = 16'sd32;
        fc1_weights[108][135] = 16'sd-8;
        fc1_weights[108][136] = 16'sd50;
        fc1_weights[108][137] = 16'sd20;
        fc1_weights[108][138] = 16'sd44;
        fc1_weights[108][139] = 16'sd40;
        fc1_weights[108][140] = 16'sd30;
        fc1_weights[108][141] = 16'sd18;
        fc1_weights[108][142] = 16'sd-10;
        fc1_weights[108][143] = 16'sd26;
        fc1_weights[108][144] = 16'sd-11;
        fc1_weights[108][145] = 16'sd15;
        fc1_weights[108][146] = 16'sd-1;
        fc1_weights[108][147] = 16'sd-32;
        fc1_weights[108][148] = 16'sd7;
        fc1_weights[108][149] = 16'sd-7;
        fc1_weights[108][150] = 16'sd-4;
        fc1_weights[108][151] = 16'sd-43;
        fc1_weights[108][152] = 16'sd-16;
        fc1_weights[108][153] = 16'sd-68;
        fc1_weights[108][154] = 16'sd2;
        fc1_weights[108][155] = 16'sd5;
        fc1_weights[108][156] = 16'sd83;
        fc1_weights[108][157] = 16'sd40;
        fc1_weights[108][158] = 16'sd31;
        fc1_weights[108][159] = 16'sd47;
        fc1_weights[108][160] = 16'sd75;
        fc1_weights[108][161] = 16'sd7;
        fc1_weights[108][162] = 16'sd31;
        fc1_weights[108][163] = 16'sd6;
        fc1_weights[108][164] = 16'sd49;
        fc1_weights[108][165] = 16'sd32;
        fc1_weights[108][166] = 16'sd49;
        fc1_weights[108][167] = 16'sd-10;
        fc1_weights[108][168] = 16'sd6;
        fc1_weights[108][169] = 16'sd-63;
        fc1_weights[108][170] = 16'sd-82;
        fc1_weights[108][171] = 16'sd-42;
        fc1_weights[108][172] = 16'sd-20;
        fc1_weights[108][173] = 16'sd-30;
        fc1_weights[108][174] = 16'sd-23;
        fc1_weights[108][175] = 16'sd-36;
        fc1_weights[108][176] = 16'sd-7;
        fc1_weights[108][177] = 16'sd-35;
        fc1_weights[108][178] = 16'sd-5;
        fc1_weights[108][179] = 16'sd-6;
        fc1_weights[108][180] = 16'sd-32;
        fc1_weights[108][181] = 16'sd27;
        fc1_weights[108][182] = 16'sd77;
        fc1_weights[108][183] = 16'sd82;
        fc1_weights[108][184] = 16'sd52;
        fc1_weights[108][185] = 16'sd-12;
        fc1_weights[108][186] = 16'sd35;
        fc1_weights[108][187] = 16'sd4;
        fc1_weights[108][188] = 16'sd37;
        fc1_weights[108][189] = 16'sd-18;
        fc1_weights[108][190] = 16'sd12;
        fc1_weights[108][191] = 16'sd4;
        fc1_weights[108][192] = 16'sd32;
        fc1_weights[108][193] = 16'sd38;
        fc1_weights[108][194] = 16'sd14;
        fc1_weights[108][195] = 16'sd-9;
        fc1_weights[108][196] = 16'sd-44;
        fc1_weights[108][197] = 16'sd-62;
        fc1_weights[108][198] = 16'sd21;
        fc1_weights[108][199] = 16'sd-4;
        fc1_weights[108][200] = 16'sd3;
        fc1_weights[108][201] = 16'sd-18;
        fc1_weights[108][202] = 16'sd-91;
        fc1_weights[108][203] = 16'sd-77;
        fc1_weights[108][204] = 16'sd-28;
        fc1_weights[108][205] = 16'sd-51;
        fc1_weights[108][206] = 16'sd-19;
        fc1_weights[108][207] = 16'sd-18;
        fc1_weights[109][0] = 16'sd-52;
        fc1_weights[109][1] = 16'sd-24;
        fc1_weights[109][2] = 16'sd1;
        fc1_weights[109][3] = 16'sd-7;
        fc1_weights[109][4] = 16'sd-24;
        fc1_weights[109][5] = 16'sd6;
        fc1_weights[109][6] = 16'sd-2;
        fc1_weights[109][7] = 16'sd-40;
        fc1_weights[109][8] = 16'sd2;
        fc1_weights[109][9] = 16'sd13;
        fc1_weights[109][10] = 16'sd-38;
        fc1_weights[109][11] = 16'sd-19;
        fc1_weights[109][12] = 16'sd56;
        fc1_weights[109][13] = 16'sd21;
        fc1_weights[109][14] = 16'sd-14;
        fc1_weights[109][15] = 16'sd-35;
        fc1_weights[109][16] = 16'sd-29;
        fc1_weights[109][17] = 16'sd29;
        fc1_weights[109][18] = 16'sd9;
        fc1_weights[109][19] = 16'sd17;
        fc1_weights[109][20] = 16'sd3;
        fc1_weights[109][21] = 16'sd20;
        fc1_weights[109][22] = 16'sd2;
        fc1_weights[109][23] = 16'sd-11;
        fc1_weights[109][24] = 16'sd-28;
        fc1_weights[109][25] = 16'sd-79;
        fc1_weights[109][26] = 16'sd-19;
        fc1_weights[109][27] = 16'sd-29;
        fc1_weights[109][28] = 16'sd-38;
        fc1_weights[109][29] = 16'sd9;
        fc1_weights[109][30] = 16'sd-9;
        fc1_weights[109][31] = 16'sd-21;
        fc1_weights[109][32] = 16'sd12;
        fc1_weights[109][33] = 16'sd-26;
        fc1_weights[109][34] = 16'sd25;
        fc1_weights[109][35] = 16'sd0;
        fc1_weights[109][36] = 16'sd-54;
        fc1_weights[109][37] = 16'sd-74;
        fc1_weights[109][38] = 16'sd-16;
        fc1_weights[109][39] = 16'sd-9;
        fc1_weights[109][40] = 16'sd-33;
        fc1_weights[109][41] = 16'sd11;
        fc1_weights[109][42] = 16'sd0;
        fc1_weights[109][43] = 16'sd-2;
        fc1_weights[109][44] = 16'sd-11;
        fc1_weights[109][45] = 16'sd79;
        fc1_weights[109][46] = 16'sd-1;
        fc1_weights[109][47] = 16'sd29;
        fc1_weights[109][48] = 16'sd25;
        fc1_weights[109][49] = 16'sd-5;
        fc1_weights[109][50] = 16'sd23;
        fc1_weights[109][51] = 16'sd39;
        fc1_weights[109][52] = 16'sd-15;
        fc1_weights[109][53] = 16'sd-21;
        fc1_weights[109][54] = 16'sd-29;
        fc1_weights[109][55] = 16'sd-14;
        fc1_weights[109][56] = 16'sd-35;
        fc1_weights[109][57] = 16'sd-73;
        fc1_weights[109][58] = 16'sd23;
        fc1_weights[109][59] = 16'sd-2;
        fc1_weights[109][60] = 16'sd-4;
        fc1_weights[109][61] = 16'sd2;
        fc1_weights[109][62] = 16'sd21;
        fc1_weights[109][63] = 16'sd-8;
        fc1_weights[109][64] = 16'sd-21;
        fc1_weights[109][65] = 16'sd9;
        fc1_weights[109][66] = 16'sd-3;
        fc1_weights[109][67] = 16'sd21;
        fc1_weights[109][68] = 16'sd15;
        fc1_weights[109][69] = 16'sd-17;
        fc1_weights[109][70] = 16'sd15;
        fc1_weights[109][71] = 16'sd-26;
        fc1_weights[109][72] = 16'sd-48;
        fc1_weights[109][73] = 16'sd26;
        fc1_weights[109][74] = 16'sd9;
        fc1_weights[109][75] = 16'sd-11;
        fc1_weights[109][76] = 16'sd1;
        fc1_weights[109][77] = 16'sd15;
        fc1_weights[109][78] = 16'sd-41;
        fc1_weights[109][79] = 16'sd-52;
        fc1_weights[109][80] = 16'sd-39;
        fc1_weights[109][81] = 16'sd1;
        fc1_weights[109][82] = 16'sd-43;
        fc1_weights[109][83] = 16'sd1;
        fc1_weights[109][84] = 16'sd11;
        fc1_weights[109][85] = 16'sd-1;
        fc1_weights[109][86] = 16'sd20;
        fc1_weights[109][87] = 16'sd21;
        fc1_weights[109][88] = 16'sd83;
        fc1_weights[109][89] = 16'sd-6;
        fc1_weights[109][90] = 16'sd-9;
        fc1_weights[109][91] = 16'sd0;
        fc1_weights[109][92] = 16'sd13;
        fc1_weights[109][93] = 16'sd-3;
        fc1_weights[109][94] = 16'sd25;
        fc1_weights[109][95] = 16'sd-27;
        fc1_weights[109][96] = 16'sd-13;
        fc1_weights[109][97] = 16'sd3;
        fc1_weights[109][98] = 16'sd24;
        fc1_weights[109][99] = 16'sd-17;
        fc1_weights[109][100] = 16'sd10;
        fc1_weights[109][101] = 16'sd-2;
        fc1_weights[109][102] = 16'sd5;
        fc1_weights[109][103] = 16'sd54;
        fc1_weights[109][104] = 16'sd-21;
        fc1_weights[109][105] = 16'sd-10;
        fc1_weights[109][106] = 16'sd-5;
        fc1_weights[109][107] = 16'sd20;
        fc1_weights[109][108] = 16'sd-7;
        fc1_weights[109][109] = 16'sd3;
        fc1_weights[109][110] = 16'sd12;
        fc1_weights[109][111] = 16'sd2;
        fc1_weights[109][112] = 16'sd-16;
        fc1_weights[109][113] = 16'sd7;
        fc1_weights[109][114] = 16'sd37;
        fc1_weights[109][115] = 16'sd33;
        fc1_weights[109][116] = 16'sd36;
        fc1_weights[109][117] = 16'sd-10;
        fc1_weights[109][118] = 16'sd-23;
        fc1_weights[109][119] = 16'sd-6;
        fc1_weights[109][120] = 16'sd18;
        fc1_weights[109][121] = 16'sd-5;
        fc1_weights[109][122] = 16'sd-47;
        fc1_weights[109][123] = 16'sd-6;
        fc1_weights[109][124] = 16'sd-3;
        fc1_weights[109][125] = 16'sd-4;
        fc1_weights[109][126] = 16'sd9;
        fc1_weights[109][127] = 16'sd10;
        fc1_weights[109][128] = 16'sd-4;
        fc1_weights[109][129] = 16'sd32;
        fc1_weights[109][130] = 16'sd-7;
        fc1_weights[109][131] = 16'sd-4;
        fc1_weights[109][132] = 16'sd-9;
        fc1_weights[109][133] = 16'sd-10;
        fc1_weights[109][134] = 16'sd-25;
        fc1_weights[109][135] = 16'sd-24;
        fc1_weights[109][136] = 16'sd-7;
        fc1_weights[109][137] = 16'sd-2;
        fc1_weights[109][138] = 16'sd-7;
        fc1_weights[109][139] = 16'sd-44;
        fc1_weights[109][140] = 16'sd-39;
        fc1_weights[109][141] = 16'sd4;
        fc1_weights[109][142] = 16'sd-26;
        fc1_weights[109][143] = 16'sd-46;
        fc1_weights[109][144] = 16'sd-3;
        fc1_weights[109][145] = 16'sd-2;
        fc1_weights[109][146] = 16'sd1;
        fc1_weights[109][147] = 16'sd-62;
        fc1_weights[109][148] = 16'sd-47;
        fc1_weights[109][149] = 16'sd-27;
        fc1_weights[109][150] = 16'sd0;
        fc1_weights[109][151] = 16'sd29;
        fc1_weights[109][152] = 16'sd-11;
        fc1_weights[109][153] = 16'sd-14;
        fc1_weights[109][154] = 16'sd41;
        fc1_weights[109][155] = 16'sd31;
        fc1_weights[109][156] = 16'sd-17;
        fc1_weights[109][157] = 16'sd-38;
        fc1_weights[109][158] = 16'sd-5;
        fc1_weights[109][159] = 16'sd41;
        fc1_weights[109][160] = 16'sd-1;
        fc1_weights[109][161] = 16'sd29;
        fc1_weights[109][162] = 16'sd39;
        fc1_weights[109][163] = 16'sd20;
        fc1_weights[109][164] = 16'sd32;
        fc1_weights[109][165] = 16'sd-3;
        fc1_weights[109][166] = 16'sd-37;
        fc1_weights[109][167] = 16'sd-44;
        fc1_weights[109][168] = 16'sd-67;
        fc1_weights[109][169] = 16'sd-35;
        fc1_weights[109][170] = 16'sd-11;
        fc1_weights[109][171] = 16'sd-48;
        fc1_weights[109][172] = 16'sd-67;
        fc1_weights[109][173] = 16'sd-73;
        fc1_weights[109][174] = 16'sd-32;
        fc1_weights[109][175] = 16'sd-14;
        fc1_weights[109][176] = 16'sd4;
        fc1_weights[109][177] = 16'sd44;
        fc1_weights[109][178] = 16'sd41;
        fc1_weights[109][179] = 16'sd43;
        fc1_weights[109][180] = 16'sd53;
        fc1_weights[109][181] = 16'sd66;
        fc1_weights[109][182] = 16'sd-3;
        fc1_weights[109][183] = 16'sd-3;
        fc1_weights[109][184] = 16'sd35;
        fc1_weights[109][185] = 16'sd4;
        fc1_weights[109][186] = 16'sd23;
        fc1_weights[109][187] = 16'sd28;
        fc1_weights[109][188] = 16'sd33;
        fc1_weights[109][189] = 16'sd44;
        fc1_weights[109][190] = 16'sd53;
        fc1_weights[109][191] = 16'sd5;
        fc1_weights[109][192] = 16'sd6;
        fc1_weights[109][193] = 16'sd-25;
        fc1_weights[109][194] = 16'sd-14;
        fc1_weights[109][195] = 16'sd5;
        fc1_weights[109][196] = 16'sd-2;
        fc1_weights[109][197] = 16'sd-6;
        fc1_weights[109][198] = 16'sd-31;
        fc1_weights[109][199] = 16'sd-14;
        fc1_weights[109][200] = 16'sd3;
        fc1_weights[109][201] = 16'sd-25;
        fc1_weights[109][202] = 16'sd26;
        fc1_weights[109][203] = 16'sd28;
        fc1_weights[109][204] = 16'sd-1;
        fc1_weights[109][205] = 16'sd42;
        fc1_weights[109][206] = 16'sd74;
        fc1_weights[109][207] = 16'sd72;
        fc1_weights[110][0] = 16'sd8;
        fc1_weights[110][1] = 16'sd10;
        fc1_weights[110][2] = 16'sd-31;
        fc1_weights[110][3] = 16'sd-13;
        fc1_weights[110][4] = 16'sd-17;
        fc1_weights[110][5] = 16'sd-16;
        fc1_weights[110][6] = 16'sd-11;
        fc1_weights[110][7] = 16'sd39;
        fc1_weights[110][8] = 16'sd-32;
        fc1_weights[110][9] = 16'sd-4;
        fc1_weights[110][10] = 16'sd-42;
        fc1_weights[110][11] = 16'sd-91;
        fc1_weights[110][12] = 16'sd-90;
        fc1_weights[110][13] = 16'sd-11;
        fc1_weights[110][14] = 16'sd24;
        fc1_weights[110][15] = 16'sd55;
        fc1_weights[110][16] = 16'sd54;
        fc1_weights[110][17] = 16'sd22;
        fc1_weights[110][18] = 16'sd-5;
        fc1_weights[110][19] = 16'sd-20;
        fc1_weights[110][20] = 16'sd46;
        fc1_weights[110][21] = 16'sd15;
        fc1_weights[110][22] = 16'sd16;
        fc1_weights[110][23] = 16'sd-57;
        fc1_weights[110][24] = 16'sd-7;
        fc1_weights[110][25] = 16'sd-13;
        fc1_weights[110][26] = 16'sd-26;
        fc1_weights[110][27] = 16'sd-19;
        fc1_weights[110][28] = 16'sd20;
        fc1_weights[110][29] = 16'sd-23;
        fc1_weights[110][30] = 16'sd-7;
        fc1_weights[110][31] = 16'sd40;
        fc1_weights[110][32] = 16'sd18;
        fc1_weights[110][33] = 16'sd-32;
        fc1_weights[110][34] = 16'sd-39;
        fc1_weights[110][35] = 16'sd-4;
        fc1_weights[110][36] = 16'sd10;
        fc1_weights[110][37] = 16'sd-78;
        fc1_weights[110][38] = 16'sd-60;
        fc1_weights[110][39] = 16'sd4;
        fc1_weights[110][40] = 16'sd57;
        fc1_weights[110][41] = 16'sd62;
        fc1_weights[110][42] = 16'sd53;
        fc1_weights[110][43] = 16'sd-60;
        fc1_weights[110][44] = 16'sd-41;
        fc1_weights[110][45] = 16'sd-95;
        fc1_weights[110][46] = 16'sd-53;
        fc1_weights[110][47] = 16'sd-9;
        fc1_weights[110][48] = 16'sd-52;
        fc1_weights[110][49] = 16'sd-43;
        fc1_weights[110][50] = 16'sd15;
        fc1_weights[110][51] = 16'sd-89;
        fc1_weights[110][52] = 16'sd-10;
        fc1_weights[110][53] = 16'sd67;
        fc1_weights[110][54] = 16'sd-18;
        fc1_weights[110][55] = 16'sd-15;
        fc1_weights[110][56] = 16'sd15;
        fc1_weights[110][57] = 16'sd14;
        fc1_weights[110][58] = 16'sd55;
        fc1_weights[110][59] = 16'sd17;
        fc1_weights[110][60] = 16'sd-31;
        fc1_weights[110][61] = 16'sd5;
        fc1_weights[110][62] = 16'sd-23;
        fc1_weights[110][63] = 16'sd27;
        fc1_weights[110][64] = 16'sd-25;
        fc1_weights[110][65] = 16'sd-29;
        fc1_weights[110][66] = 16'sd37;
        fc1_weights[110][67] = 16'sd15;
        fc1_weights[110][68] = 16'sd9;
        fc1_weights[110][69] = 16'sd-52;
        fc1_weights[110][70] = 16'sd-79;
        fc1_weights[110][71] = 16'sd-35;
        fc1_weights[110][72] = 16'sd30;
        fc1_weights[110][73] = 16'sd-23;
        fc1_weights[110][74] = 16'sd-22;
        fc1_weights[110][75] = 16'sd-26;
        fc1_weights[110][76] = 16'sd-67;
        fc1_weights[110][77] = 16'sd-34;
        fc1_weights[110][78] = 16'sd29;
        fc1_weights[110][79] = 16'sd115;
        fc1_weights[110][80] = 16'sd22;
        fc1_weights[110][81] = 16'sd0;
        fc1_weights[110][82] = 16'sd32;
        fc1_weights[110][83] = 16'sd48;
        fc1_weights[110][84] = 16'sd49;
        fc1_weights[110][85] = 16'sd17;
        fc1_weights[110][86] = 16'sd48;
        fc1_weights[110][87] = 16'sd-57;
        fc1_weights[110][88] = 16'sd-49;
        fc1_weights[110][89] = 16'sd-60;
        fc1_weights[110][90] = 16'sd9;
        fc1_weights[110][91] = 16'sd29;
        fc1_weights[110][92] = 16'sd31;
        fc1_weights[110][93] = 16'sd47;
        fc1_weights[110][94] = 16'sd12;
        fc1_weights[110][95] = 16'sd31;
        fc1_weights[110][96] = 16'sd-28;
        fc1_weights[110][97] = 16'sd-11;
        fc1_weights[110][98] = 16'sd46;
        fc1_weights[110][99] = 16'sd51;
        fc1_weights[110][100] = 16'sd9;
        fc1_weights[110][101] = 16'sd-7;
        fc1_weights[110][102] = 16'sd0;
        fc1_weights[110][103] = 16'sd-43;
        fc1_weights[110][104] = 16'sd29;
        fc1_weights[110][105] = 16'sd-6;
        fc1_weights[110][106] = 16'sd40;
        fc1_weights[110][107] = 16'sd4;
        fc1_weights[110][108] = 16'sd52;
        fc1_weights[110][109] = 16'sd6;
        fc1_weights[110][110] = 16'sd37;
        fc1_weights[110][111] = 16'sd-23;
        fc1_weights[110][112] = 16'sd8;
        fc1_weights[110][113] = 16'sd-3;
        fc1_weights[110][114] = 16'sd-46;
        fc1_weights[110][115] = 16'sd-24;
        fc1_weights[110][116] = 16'sd-72;
        fc1_weights[110][117] = 16'sd-7;
        fc1_weights[110][118] = 16'sd10;
        fc1_weights[110][119] = 16'sd23;
        fc1_weights[110][120] = 16'sd23;
        fc1_weights[110][121] = 16'sd-8;
        fc1_weights[110][122] = 16'sd-18;
        fc1_weights[110][123] = 16'sd-4;
        fc1_weights[110][124] = 16'sd3;
        fc1_weights[110][125] = 16'sd4;
        fc1_weights[110][126] = 16'sd-66;
        fc1_weights[110][127] = 16'sd-6;
        fc1_weights[110][128] = 16'sd-20;
        fc1_weights[110][129] = 16'sd-127;
        fc1_weights[110][130] = 16'sd-53;
        fc1_weights[110][131] = 16'sd-27;
        fc1_weights[110][132] = 16'sd-10;
        fc1_weights[110][133] = 16'sd-49;
        fc1_weights[110][134] = 16'sd-12;
        fc1_weights[110][135] = 16'sd-18;
        fc1_weights[110][136] = 16'sd-9;
        fc1_weights[110][137] = 16'sd53;
        fc1_weights[110][138] = 16'sd5;
        fc1_weights[110][139] = 16'sd30;
        fc1_weights[110][140] = 16'sd70;
        fc1_weights[110][141] = 16'sd54;
        fc1_weights[110][142] = 16'sd39;
        fc1_weights[110][143] = 16'sd-3;
        fc1_weights[110][144] = 16'sd0;
        fc1_weights[110][145] = 16'sd-23;
        fc1_weights[110][146] = 16'sd-49;
        fc1_weights[110][147] = 16'sd41;
        fc1_weights[110][148] = 16'sd-10;
        fc1_weights[110][149] = 16'sd-65;
        fc1_weights[110][150] = 16'sd-49;
        fc1_weights[110][151] = 16'sd-9;
        fc1_weights[110][152] = 16'sd-11;
        fc1_weights[110][153] = 16'sd12;
        fc1_weights[110][154] = 16'sd0;
        fc1_weights[110][155] = 16'sd7;
        fc1_weights[110][156] = 16'sd-28;
        fc1_weights[110][157] = 16'sd51;
        fc1_weights[110][158] = 16'sd0;
        fc1_weights[110][159] = 16'sd-40;
        fc1_weights[110][160] = 16'sd-29;
        fc1_weights[110][161] = 16'sd-24;
        fc1_weights[110][162] = 16'sd-39;
        fc1_weights[110][163] = 16'sd22;
        fc1_weights[110][164] = 16'sd-15;
        fc1_weights[110][165] = 16'sd-2;
        fc1_weights[110][166] = 16'sd18;
        fc1_weights[110][167] = 16'sd57;
        fc1_weights[110][168] = 16'sd-8;
        fc1_weights[110][169] = 16'sd6;
        fc1_weights[110][170] = 16'sd12;
        fc1_weights[110][171] = 16'sd8;
        fc1_weights[110][172] = 16'sd10;
        fc1_weights[110][173] = 16'sd25;
        fc1_weights[110][174] = 16'sd-3;
        fc1_weights[110][175] = 16'sd22;
        fc1_weights[110][176] = 16'sd-9;
        fc1_weights[110][177] = 16'sd10;
        fc1_weights[110][178] = 16'sd-1;
        fc1_weights[110][179] = 16'sd-7;
        fc1_weights[110][180] = 16'sd6;
        fc1_weights[110][181] = 16'sd-16;
        fc1_weights[110][182] = 16'sd-6;
        fc1_weights[110][183] = 16'sd-11;
        fc1_weights[110][184] = 16'sd-42;
        fc1_weights[110][185] = 16'sd-11;
        fc1_weights[110][186] = 16'sd7;
        fc1_weights[110][187] = 16'sd7;
        fc1_weights[110][188] = 16'sd-43;
        fc1_weights[110][189] = 16'sd9;
        fc1_weights[110][190] = 16'sd12;
        fc1_weights[110][191] = 16'sd11;
        fc1_weights[110][192] = 16'sd23;
        fc1_weights[110][193] = 16'sd22;
        fc1_weights[110][194] = 16'sd49;
        fc1_weights[110][195] = 16'sd63;
        fc1_weights[110][196] = 16'sd27;
        fc1_weights[110][197] = 16'sd4;
        fc1_weights[110][198] = 16'sd-31;
        fc1_weights[110][199] = 16'sd84;
        fc1_weights[110][200] = 16'sd-15;
        fc1_weights[110][201] = 16'sd-46;
        fc1_weights[110][202] = 16'sd25;
        fc1_weights[110][203] = 16'sd18;
        fc1_weights[110][204] = 16'sd-17;
        fc1_weights[110][205] = 16'sd10;
        fc1_weights[110][206] = 16'sd-26;
        fc1_weights[110][207] = 16'sd-16;
        fc1_weights[111][0] = 16'sd5;
        fc1_weights[111][1] = 16'sd28;
        fc1_weights[111][2] = 16'sd0;
        fc1_weights[111][3] = 16'sd3;
        fc1_weights[111][4] = 16'sd-16;
        fc1_weights[111][5] = 16'sd-13;
        fc1_weights[111][6] = 16'sd-1;
        fc1_weights[111][7] = 16'sd-8;
        fc1_weights[111][8] = 16'sd-25;
        fc1_weights[111][9] = 16'sd-73;
        fc1_weights[111][10] = 16'sd-29;
        fc1_weights[111][11] = 16'sd-51;
        fc1_weights[111][12] = 16'sd-43;
        fc1_weights[111][13] = 16'sd-5;
        fc1_weights[111][14] = 16'sd-1;
        fc1_weights[111][15] = 16'sd37;
        fc1_weights[111][16] = 16'sd35;
        fc1_weights[111][17] = 16'sd42;
        fc1_weights[111][18] = 16'sd16;
        fc1_weights[111][19] = 16'sd-35;
        fc1_weights[111][20] = 16'sd-28;
        fc1_weights[111][21] = 16'sd-23;
        fc1_weights[111][22] = 16'sd-41;
        fc1_weights[111][23] = 16'sd-27;
        fc1_weights[111][24] = 16'sd-9;
        fc1_weights[111][25] = 16'sd-8;
        fc1_weights[111][26] = 16'sd10;
        fc1_weights[111][27] = 16'sd1;
        fc1_weights[111][28] = 16'sd8;
        fc1_weights[111][29] = 16'sd6;
        fc1_weights[111][30] = 16'sd-6;
        fc1_weights[111][31] = 16'sd29;
        fc1_weights[111][32] = 16'sd-11;
        fc1_weights[111][33] = 16'sd-38;
        fc1_weights[111][34] = 16'sd-26;
        fc1_weights[111][35] = 16'sd-40;
        fc1_weights[111][36] = 16'sd-12;
        fc1_weights[111][37] = 16'sd-47;
        fc1_weights[111][38] = 16'sd-50;
        fc1_weights[111][39] = 16'sd-27;
        fc1_weights[111][40] = 16'sd-10;
        fc1_weights[111][41] = 16'sd19;
        fc1_weights[111][42] = 16'sd30;
        fc1_weights[111][43] = 16'sd-20;
        fc1_weights[111][44] = 16'sd-10;
        fc1_weights[111][45] = 16'sd-44;
        fc1_weights[111][46] = 16'sd-62;
        fc1_weights[111][47] = 16'sd-50;
        fc1_weights[111][48] = 16'sd-22;
        fc1_weights[111][49] = 16'sd-26;
        fc1_weights[111][50] = 16'sd-6;
        fc1_weights[111][51] = 16'sd-11;
        fc1_weights[111][52] = 16'sd35;
        fc1_weights[111][53] = 16'sd52;
        fc1_weights[111][54] = 16'sd-5;
        fc1_weights[111][55] = 16'sd13;
        fc1_weights[111][56] = 16'sd33;
        fc1_weights[111][57] = 16'sd40;
        fc1_weights[111][58] = 16'sd32;
        fc1_weights[111][59] = 16'sd-7;
        fc1_weights[111][60] = 16'sd-20;
        fc1_weights[111][61] = 16'sd-6;
        fc1_weights[111][62] = 16'sd-30;
        fc1_weights[111][63] = 16'sd-22;
        fc1_weights[111][64] = 16'sd-25;
        fc1_weights[111][65] = 16'sd-37;
        fc1_weights[111][66] = 16'sd24;
        fc1_weights[111][67] = 16'sd-7;
        fc1_weights[111][68] = 16'sd-11;
        fc1_weights[111][69] = 16'sd-5;
        fc1_weights[111][70] = 16'sd38;
        fc1_weights[111][71] = 16'sd-14;
        fc1_weights[111][72] = 16'sd-39;
        fc1_weights[111][73] = 16'sd-19;
        fc1_weights[111][74] = 16'sd-4;
        fc1_weights[111][75] = 16'sd-2;
        fc1_weights[111][76] = 16'sd15;
        fc1_weights[111][77] = 16'sd-5;
        fc1_weights[111][78] = 16'sd9;
        fc1_weights[111][79] = 16'sd23;
        fc1_weights[111][80] = 16'sd-2;
        fc1_weights[111][81] = 16'sd35;
        fc1_weights[111][82] = 16'sd-4;
        fc1_weights[111][83] = 16'sd43;
        fc1_weights[111][84] = 16'sd-4;
        fc1_weights[111][85] = 16'sd5;
        fc1_weights[111][86] = 16'sd18;
        fc1_weights[111][87] = 16'sd21;
        fc1_weights[111][88] = 16'sd55;
        fc1_weights[111][89] = 16'sd0;
        fc1_weights[111][90] = 16'sd-8;
        fc1_weights[111][91] = 16'sd5;
        fc1_weights[111][92] = 16'sd28;
        fc1_weights[111][93] = 16'sd23;
        fc1_weights[111][94] = 16'sd-36;
        fc1_weights[111][95] = 16'sd5;
        fc1_weights[111][96] = 16'sd0;
        fc1_weights[111][97] = 16'sd5;
        fc1_weights[111][98] = 16'sd8;
        fc1_weights[111][99] = 16'sd-8;
        fc1_weights[111][100] = 16'sd4;
        fc1_weights[111][101] = 16'sd-24;
        fc1_weights[111][102] = 16'sd4;
        fc1_weights[111][103] = 16'sd-7;
        fc1_weights[111][104] = 16'sd17;
        fc1_weights[111][105] = 16'sd-19;
        fc1_weights[111][106] = 16'sd41;
        fc1_weights[111][107] = 16'sd52;
        fc1_weights[111][108] = 16'sd36;
        fc1_weights[111][109] = 16'sd11;
        fc1_weights[111][110] = 16'sd-3;
        fc1_weights[111][111] = 16'sd-8;
        fc1_weights[111][112] = 16'sd32;
        fc1_weights[111][113] = 16'sd27;
        fc1_weights[111][114] = 16'sd-14;
        fc1_weights[111][115] = 16'sd-6;
        fc1_weights[111][116] = 16'sd-24;
        fc1_weights[111][117] = 16'sd8;
        fc1_weights[111][118] = 16'sd-13;
        fc1_weights[111][119] = 16'sd-14;
        fc1_weights[111][120] = 16'sd-8;
        fc1_weights[111][121] = 16'sd-16;
        fc1_weights[111][122] = 16'sd-3;
        fc1_weights[111][123] = 16'sd-4;
        fc1_weights[111][124] = 16'sd-30;
        fc1_weights[111][125] = 16'sd-40;
        fc1_weights[111][126] = 16'sd-33;
        fc1_weights[111][127] = 16'sd-15;
        fc1_weights[111][128] = 16'sd5;
        fc1_weights[111][129] = 16'sd-11;
        fc1_weights[111][130] = 16'sd-7;
        fc1_weights[111][131] = 16'sd4;
        fc1_weights[111][132] = 16'sd6;
        fc1_weights[111][133] = 16'sd12;
        fc1_weights[111][134] = 16'sd-11;
        fc1_weights[111][135] = 16'sd-1;
        fc1_weights[111][136] = 16'sd-4;
        fc1_weights[111][137] = 16'sd2;
        fc1_weights[111][138] = 16'sd-38;
        fc1_weights[111][139] = 16'sd-24;
        fc1_weights[111][140] = 16'sd1;
        fc1_weights[111][141] = 16'sd23;
        fc1_weights[111][142] = 16'sd39;
        fc1_weights[111][143] = 16'sd2;
        fc1_weights[111][144] = 16'sd18;
        fc1_weights[111][145] = 16'sd-6;
        fc1_weights[111][146] = 16'sd-16;
        fc1_weights[111][147] = 16'sd-7;
        fc1_weights[111][148] = 16'sd-16;
        fc1_weights[111][149] = 16'sd-36;
        fc1_weights[111][150] = 16'sd-27;
        fc1_weights[111][151] = 16'sd-30;
        fc1_weights[111][152] = 16'sd2;
        fc1_weights[111][153] = 16'sd-2;
        fc1_weights[111][154] = 16'sd8;
        fc1_weights[111][155] = 16'sd-14;
        fc1_weights[111][156] = 16'sd14;
        fc1_weights[111][157] = 16'sd49;
        fc1_weights[111][158] = 16'sd10;
        fc1_weights[111][159] = 16'sd8;
        fc1_weights[111][160] = 16'sd17;
        fc1_weights[111][161] = 16'sd-9;
        fc1_weights[111][162] = 16'sd12;
        fc1_weights[111][163] = 16'sd32;
        fc1_weights[111][164] = 16'sd-2;
        fc1_weights[111][165] = 16'sd14;
        fc1_weights[111][166] = 16'sd-28;
        fc1_weights[111][167] = 16'sd-21;
        fc1_weights[111][168] = 16'sd-30;
        fc1_weights[111][169] = 16'sd-6;
        fc1_weights[111][170] = 16'sd-26;
        fc1_weights[111][171] = 16'sd-11;
        fc1_weights[111][172] = 16'sd-30;
        fc1_weights[111][173] = 16'sd1;
        fc1_weights[111][174] = 16'sd-24;
        fc1_weights[111][175] = 16'sd-3;
        fc1_weights[111][176] = 16'sd-20;
        fc1_weights[111][177] = 16'sd-12;
        fc1_weights[111][178] = 16'sd-12;
        fc1_weights[111][179] = 16'sd-26;
        fc1_weights[111][180] = 16'sd4;
        fc1_weights[111][181] = 16'sd-8;
        fc1_weights[111][182] = 16'sd13;
        fc1_weights[111][183] = 16'sd20;
        fc1_weights[111][184] = 16'sd-4;
        fc1_weights[111][185] = 16'sd21;
        fc1_weights[111][186] = 16'sd2;
        fc1_weights[111][187] = 16'sd-22;
        fc1_weights[111][188] = 16'sd-26;
        fc1_weights[111][189] = 16'sd14;
        fc1_weights[111][190] = 16'sd8;
        fc1_weights[111][191] = 16'sd-10;
        fc1_weights[111][192] = 16'sd-1;
        fc1_weights[111][193] = 16'sd-26;
        fc1_weights[111][194] = 16'sd1;
        fc1_weights[111][195] = 16'sd6;
        fc1_weights[111][196] = 16'sd-14;
        fc1_weights[111][197] = 16'sd3;
        fc1_weights[111][198] = 16'sd-1;
        fc1_weights[111][199] = 16'sd45;
        fc1_weights[111][200] = 16'sd-7;
        fc1_weights[111][201] = 16'sd2;
        fc1_weights[111][202] = 16'sd-3;
        fc1_weights[111][203] = 16'sd20;
        fc1_weights[111][204] = 16'sd1;
        fc1_weights[111][205] = 16'sd-4;
        fc1_weights[111][206] = 16'sd-35;
        fc1_weights[111][207] = 16'sd-7;
        fc1_weights[112][0] = 16'sd-13;
        fc1_weights[112][1] = 16'sd-123;
        fc1_weights[112][2] = 16'sd-56;
        fc1_weights[112][3] = 16'sd-22;
        fc1_weights[112][4] = 16'sd-35;
        fc1_weights[112][5] = 16'sd-21;
        fc1_weights[112][6] = 16'sd12;
        fc1_weights[112][7] = 16'sd2;
        fc1_weights[112][8] = 16'sd29;
        fc1_weights[112][9] = 16'sd-76;
        fc1_weights[112][10] = 16'sd-9;
        fc1_weights[112][11] = 16'sd61;
        fc1_weights[112][12] = 16'sd171;
        fc1_weights[112][13] = 16'sd54;
        fc1_weights[112][14] = 16'sd78;
        fc1_weights[112][15] = 16'sd-18;
        fc1_weights[112][16] = 16'sd-41;
        fc1_weights[112][17] = 16'sd-3;
        fc1_weights[112][18] = 16'sd38;
        fc1_weights[112][19] = 16'sd84;
        fc1_weights[112][20] = 16'sd-16;
        fc1_weights[112][21] = 16'sd25;
        fc1_weights[112][22] = 16'sd11;
        fc1_weights[112][23] = 16'sd11;
        fc1_weights[112][24] = 16'sd-31;
        fc1_weights[112][25] = 16'sd-46;
        fc1_weights[112][26] = 16'sd5;
        fc1_weights[112][27] = 16'sd-26;
        fc1_weights[112][28] = 16'sd-34;
        fc1_weights[112][29] = 16'sd-5;
        fc1_weights[112][30] = 16'sd-27;
        fc1_weights[112][31] = 16'sd-13;
        fc1_weights[112][32] = 16'sd14;
        fc1_weights[112][33] = 16'sd78;
        fc1_weights[112][34] = 16'sd46;
        fc1_weights[112][35] = 16'sd-1;
        fc1_weights[112][36] = 16'sd-56;
        fc1_weights[112][37] = 16'sd16;
        fc1_weights[112][38] = 16'sd67;
        fc1_weights[112][39] = 16'sd44;
        fc1_weights[112][40] = 16'sd-17;
        fc1_weights[112][41] = 16'sd9;
        fc1_weights[112][42] = 16'sd45;
        fc1_weights[112][43] = 16'sd-11;
        fc1_weights[112][44] = 16'sd-4;
        fc1_weights[112][45] = 16'sd59;
        fc1_weights[112][46] = 16'sd80;
        fc1_weights[112][47] = 16'sd-8;
        fc1_weights[112][48] = 16'sd11;
        fc1_weights[112][49] = 16'sd-14;
        fc1_weights[112][50] = 16'sd-10;
        fc1_weights[112][51] = 16'sd39;
        fc1_weights[112][52] = 16'sd37;
        fc1_weights[112][53] = 16'sd-1;
        fc1_weights[112][54] = 16'sd29;
        fc1_weights[112][55] = 16'sd4;
        fc1_weights[112][56] = 16'sd-17;
        fc1_weights[112][57] = 16'sd-39;
        fc1_weights[112][58] = 16'sd-6;
        fc1_weights[112][59] = 16'sd-9;
        fc1_weights[112][60] = 16'sd-26;
        fc1_weights[112][61] = 16'sd-77;
        fc1_weights[112][62] = 16'sd43;
        fc1_weights[112][63] = 16'sd-3;
        fc1_weights[112][64] = 16'sd5;
        fc1_weights[112][65] = 16'sd74;
        fc1_weights[112][66] = 16'sd-49;
        fc1_weights[112][67] = 16'sd-35;
        fc1_weights[112][68] = 16'sd-41;
        fc1_weights[112][69] = 16'sd15;
        fc1_weights[112][70] = 16'sd7;
        fc1_weights[112][71] = 16'sd64;
        fc1_weights[112][72] = 16'sd-21;
        fc1_weights[112][73] = 16'sd-7;
        fc1_weights[112][74] = 16'sd-22;
        fc1_weights[112][75] = 16'sd7;
        fc1_weights[112][76] = 16'sd3;
        fc1_weights[112][77] = 16'sd31;
        fc1_weights[112][78] = 16'sd45;
        fc1_weights[112][79] = 16'sd-24;
        fc1_weights[112][80] = 16'sd-14;
        fc1_weights[112][81] = 16'sd13;
        fc1_weights[112][82] = 16'sd16;
        fc1_weights[112][83] = 16'sd20;
        fc1_weights[112][84] = 16'sd18;
        fc1_weights[112][85] = 16'sd0;
        fc1_weights[112][86] = 16'sd-47;
        fc1_weights[112][87] = 16'sd2;
        fc1_weights[112][88] = 16'sd35;
        fc1_weights[112][89] = 16'sd34;
        fc1_weights[112][90] = 16'sd-14;
        fc1_weights[112][91] = 16'sd-65;
        fc1_weights[112][92] = 16'sd-9;
        fc1_weights[112][93] = 16'sd-129;
        fc1_weights[112][94] = 16'sd-77;
        fc1_weights[112][95] = 16'sd-44;
        fc1_weights[112][96] = 16'sd-10;
        fc1_weights[112][97] = 16'sd11;
        fc1_weights[112][98] = 16'sd-33;
        fc1_weights[112][99] = 16'sd-15;
        fc1_weights[112][100] = 16'sd-32;
        fc1_weights[112][101] = 16'sd7;
        fc1_weights[112][102] = 16'sd-2;
        fc1_weights[112][103] = 16'sd39;
        fc1_weights[112][104] = 16'sd42;
        fc1_weights[112][105] = 16'sd49;
        fc1_weights[112][106] = 16'sd-51;
        fc1_weights[112][107] = 16'sd-25;
        fc1_weights[112][108] = 16'sd-11;
        fc1_weights[112][109] = 16'sd-9;
        fc1_weights[112][110] = 16'sd-30;
        fc1_weights[112][111] = 16'sd-34;
        fc1_weights[112][112] = 16'sd-120;
        fc1_weights[112][113] = 16'sd-11;
        fc1_weights[112][114] = 16'sd7;
        fc1_weights[112][115] = 16'sd4;
        fc1_weights[112][116] = 16'sd-17;
        fc1_weights[112][117] = 16'sd-32;
        fc1_weights[112][118] = 16'sd-23;
        fc1_weights[112][119] = 16'sd-40;
        fc1_weights[112][120] = 16'sd-11;
        fc1_weights[112][121] = 16'sd-63;
        fc1_weights[112][122] = 16'sd-101;
        fc1_weights[112][123] = 16'sd-21;
        fc1_weights[112][124] = 16'sd59;
        fc1_weights[112][125] = 16'sd-30;
        fc1_weights[112][126] = 16'sd82;
        fc1_weights[112][127] = 16'sd-17;
        fc1_weights[112][128] = 16'sd51;
        fc1_weights[112][129] = 16'sd75;
        fc1_weights[112][130] = 16'sd51;
        fc1_weights[112][131] = 16'sd5;
        fc1_weights[112][132] = 16'sd4;
        fc1_weights[112][133] = 16'sd17;
        fc1_weights[112][134] = 16'sd-31;
        fc1_weights[112][135] = 16'sd-8;
        fc1_weights[112][136] = 16'sd-25;
        fc1_weights[112][137] = 16'sd13;
        fc1_weights[112][138] = 16'sd-53;
        fc1_weights[112][139] = 16'sd-31;
        fc1_weights[112][140] = 16'sd-28;
        fc1_weights[112][141] = 16'sd-5;
        fc1_weights[112][142] = 16'sd-60;
        fc1_weights[112][143] = 16'sd11;
        fc1_weights[112][144] = 16'sd38;
        fc1_weights[112][145] = 16'sd41;
        fc1_weights[112][146] = 16'sd20;
        fc1_weights[112][147] = 16'sd0;
        fc1_weights[112][148] = 16'sd-14;
        fc1_weights[112][149] = 16'sd-4;
        fc1_weights[112][150] = 16'sd9;
        fc1_weights[112][151] = 16'sd-27;
        fc1_weights[112][152] = 16'sd-1;
        fc1_weights[112][153] = 16'sd-82;
        fc1_weights[112][154] = 16'sd-16;
        fc1_weights[112][155] = 16'sd-77;
        fc1_weights[112][156] = 16'sd17;
        fc1_weights[112][157] = 16'sd-23;
        fc1_weights[112][158] = 16'sd63;
        fc1_weights[112][159] = 16'sd90;
        fc1_weights[112][160] = 16'sd-5;
        fc1_weights[112][161] = 16'sd-20;
        fc1_weights[112][162] = 16'sd-25;
        fc1_weights[112][163] = 16'sd-13;
        fc1_weights[112][164] = 16'sd41;
        fc1_weights[112][165] = 16'sd100;
        fc1_weights[112][166] = 16'sd29;
        fc1_weights[112][167] = 16'sd10;
        fc1_weights[112][168] = 16'sd17;
        fc1_weights[112][169] = 16'sd11;
        fc1_weights[112][170] = 16'sd-26;
        fc1_weights[112][171] = 16'sd48;
        fc1_weights[112][172] = 16'sd-35;
        fc1_weights[112][173] = 16'sd-12;
        fc1_weights[112][174] = 16'sd0;
        fc1_weights[112][175] = 16'sd15;
        fc1_weights[112][176] = 16'sd-43;
        fc1_weights[112][177] = 16'sd-82;
        fc1_weights[112][178] = 16'sd15;
        fc1_weights[112][179] = 16'sd-88;
        fc1_weights[112][180] = 16'sd-74;
        fc1_weights[112][181] = 16'sd-61;
        fc1_weights[112][182] = 16'sd16;
        fc1_weights[112][183] = 16'sd7;
        fc1_weights[112][184] = 16'sd-30;
        fc1_weights[112][185] = 16'sd-27;
        fc1_weights[112][186] = 16'sd14;
        fc1_weights[112][187] = 16'sd-26;
        fc1_weights[112][188] = 16'sd15;
        fc1_weights[112][189] = 16'sd20;
        fc1_weights[112][190] = 16'sd14;
        fc1_weights[112][191] = 16'sd-55;
        fc1_weights[112][192] = 16'sd15;
        fc1_weights[112][193] = 16'sd44;
        fc1_weights[112][194] = 16'sd32;
        fc1_weights[112][195] = 16'sd42;
        fc1_weights[112][196] = 16'sd66;
        fc1_weights[112][197] = 16'sd-40;
        fc1_weights[112][198] = 16'sd61;
        fc1_weights[112][199] = 16'sd-56;
        fc1_weights[112][200] = 16'sd-22;
        fc1_weights[112][201] = 16'sd24;
        fc1_weights[112][202] = 16'sd-30;
        fc1_weights[112][203] = 16'sd-35;
        fc1_weights[112][204] = 16'sd-67;
        fc1_weights[112][205] = 16'sd-47;
        fc1_weights[112][206] = 16'sd-15;
        fc1_weights[112][207] = 16'sd-20;
        fc1_weights[113][0] = 16'sd44;
        fc1_weights[113][1] = 16'sd11;
        fc1_weights[113][2] = 16'sd11;
        fc1_weights[113][3] = 16'sd18;
        fc1_weights[113][4] = 16'sd17;
        fc1_weights[113][5] = 16'sd-24;
        fc1_weights[113][6] = 16'sd11;
        fc1_weights[113][7] = 16'sd-24;
        fc1_weights[113][8] = 16'sd-11;
        fc1_weights[113][9] = 16'sd-23;
        fc1_weights[113][10] = 16'sd-44;
        fc1_weights[113][11] = 16'sd107;
        fc1_weights[113][12] = 16'sd98;
        fc1_weights[113][13] = 16'sd72;
        fc1_weights[113][14] = 16'sd0;
        fc1_weights[113][15] = 16'sd-50;
        fc1_weights[113][16] = 16'sd-46;
        fc1_weights[113][17] = 16'sd-7;
        fc1_weights[113][18] = 16'sd-47;
        fc1_weights[113][19] = 16'sd46;
        fc1_weights[113][20] = 16'sd44;
        fc1_weights[113][21] = 16'sd24;
        fc1_weights[113][22] = 16'sd23;
        fc1_weights[113][23] = 16'sd69;
        fc1_weights[113][24] = 16'sd-9;
        fc1_weights[113][25] = 16'sd-69;
        fc1_weights[113][26] = 16'sd11;
        fc1_weights[113][27] = 16'sd43;
        fc1_weights[113][28] = 16'sd-6;
        fc1_weights[113][29] = 16'sd12;
        fc1_weights[113][30] = 16'sd-52;
        fc1_weights[113][31] = 16'sd-6;
        fc1_weights[113][32] = 16'sd36;
        fc1_weights[113][33] = 16'sd74;
        fc1_weights[113][34] = 16'sd51;
        fc1_weights[113][35] = 16'sd6;
        fc1_weights[113][36] = 16'sd-36;
        fc1_weights[113][37] = 16'sd-20;
        fc1_weights[113][38] = 16'sd121;
        fc1_weights[113][39] = 16'sd92;
        fc1_weights[113][40] = 16'sd-37;
        fc1_weights[113][41] = 16'sd-3;
        fc1_weights[113][42] = 16'sd32;
        fc1_weights[113][43] = 16'sd-21;
        fc1_weights[113][44] = 16'sd52;
        fc1_weights[113][45] = 16'sd71;
        fc1_weights[113][46] = 16'sd13;
        fc1_weights[113][47] = 16'sd35;
        fc1_weights[113][48] = 16'sd43;
        fc1_weights[113][49] = 16'sd0;
        fc1_weights[113][50] = 16'sd-17;
        fc1_weights[113][51] = 16'sd41;
        fc1_weights[113][52] = 16'sd17;
        fc1_weights[113][53] = 16'sd17;
        fc1_weights[113][54] = 16'sd36;
        fc1_weights[113][55] = 16'sd-43;
        fc1_weights[113][56] = 16'sd45;
        fc1_weights[113][57] = 16'sd-32;
        fc1_weights[113][58] = 16'sd23;
        fc1_weights[113][59] = 16'sd64;
        fc1_weights[113][60] = 16'sd15;
        fc1_weights[113][61] = 16'sd6;
        fc1_weights[113][62] = 16'sd77;
        fc1_weights[113][63] = 16'sd-15;
        fc1_weights[113][64] = 16'sd16;
        fc1_weights[113][65] = 16'sd61;
        fc1_weights[113][66] = 16'sd-17;
        fc1_weights[113][67] = 16'sd-58;
        fc1_weights[113][68] = 16'sd-13;
        fc1_weights[113][69] = 16'sd-45;
        fc1_weights[113][70] = 16'sd-48;
        fc1_weights[113][71] = 16'sd5;
        fc1_weights[113][72] = 16'sd14;
        fc1_weights[113][73] = 16'sd-39;
        fc1_weights[113][74] = 16'sd-30;
        fc1_weights[113][75] = 16'sd-5;
        fc1_weights[113][76] = 16'sd-32;
        fc1_weights[113][77] = 16'sd-18;
        fc1_weights[113][78] = 16'sd-53;
        fc1_weights[113][79] = 16'sd-101;
        fc1_weights[113][80] = 16'sd-19;
        fc1_weights[113][81] = 16'sd-54;
        fc1_weights[113][82] = 16'sd33;
        fc1_weights[113][83] = 16'sd16;
        fc1_weights[113][84] = 16'sd31;
        fc1_weights[113][85] = 16'sd45;
        fc1_weights[113][86] = 16'sd4;
        fc1_weights[113][87] = 16'sd-66;
        fc1_weights[113][88] = 16'sd-47;
        fc1_weights[113][89] = 16'sd-11;
        fc1_weights[113][90] = 16'sd48;
        fc1_weights[113][91] = 16'sd2;
        fc1_weights[113][92] = 16'sd6;
        fc1_weights[113][93] = 16'sd-82;
        fc1_weights[113][94] = 16'sd-31;
        fc1_weights[113][95] = 16'sd-67;
        fc1_weights[113][96] = 16'sd-20;
        fc1_weights[113][97] = 16'sd-27;
        fc1_weights[113][98] = 16'sd11;
        fc1_weights[113][99] = 16'sd-10;
        fc1_weights[113][100] = 16'sd29;
        fc1_weights[113][101] = 16'sd20;
        fc1_weights[113][102] = 16'sd-20;
        fc1_weights[113][103] = 16'sd43;
        fc1_weights[113][104] = 16'sd-24;
        fc1_weights[113][105] = 16'sd14;
        fc1_weights[113][106] = 16'sd-21;
        fc1_weights[113][107] = 16'sd-28;
        fc1_weights[113][108] = 16'sd-8;
        fc1_weights[113][109] = 16'sd-38;
        fc1_weights[113][110] = 16'sd3;
        fc1_weights[113][111] = 16'sd15;
        fc1_weights[113][112] = 16'sd-117;
        fc1_weights[113][113] = 16'sd-1;
        fc1_weights[113][114] = 16'sd45;
        fc1_weights[113][115] = 16'sd106;
        fc1_weights[113][116] = 16'sd-19;
        fc1_weights[113][117] = 16'sd-103;
        fc1_weights[113][118] = 16'sd-3;
        fc1_weights[113][119] = 16'sd-56;
        fc1_weights[113][120] = 16'sd-90;
        fc1_weights[113][121] = 16'sd-24;
        fc1_weights[113][122] = 16'sd-57;
        fc1_weights[113][123] = 16'sd-104;
        fc1_weights[113][124] = 16'sd-9;
        fc1_weights[113][125] = 16'sd-45;
        fc1_weights[113][126] = 16'sd72;
        fc1_weights[113][127] = 16'sd-44;
        fc1_weights[113][128] = 16'sd33;
        fc1_weights[113][129] = 16'sd60;
        fc1_weights[113][130] = 16'sd45;
        fc1_weights[113][131] = 16'sd57;
        fc1_weights[113][132] = 16'sd0;
        fc1_weights[113][133] = 16'sd20;
        fc1_weights[113][134] = 16'sd71;
        fc1_weights[113][135] = 16'sd57;
        fc1_weights[113][136] = 16'sd37;
        fc1_weights[113][137] = 16'sd57;
        fc1_weights[113][138] = 16'sd21;
        fc1_weights[113][139] = 16'sd63;
        fc1_weights[113][140] = 16'sd13;
        fc1_weights[113][141] = 16'sd62;
        fc1_weights[113][142] = 16'sd-2;
        fc1_weights[113][143] = 16'sd80;
        fc1_weights[113][144] = 16'sd-6;
        fc1_weights[113][145] = 16'sd87;
        fc1_weights[113][146] = 16'sd53;
        fc1_weights[113][147] = 16'sd-22;
        fc1_weights[113][148] = 16'sd-23;
        fc1_weights[113][149] = 16'sd33;
        fc1_weights[113][150] = 16'sd0;
        fc1_weights[113][151] = 16'sd-32;
        fc1_weights[113][152] = 16'sd6;
        fc1_weights[113][153] = 16'sd-37;
        fc1_weights[113][154] = 16'sd4;
        fc1_weights[113][155] = 16'sd-34;
        fc1_weights[113][156] = 16'sd-12;
        fc1_weights[113][157] = 16'sd-33;
        fc1_weights[113][158] = 16'sd53;
        fc1_weights[113][159] = 16'sd27;
        fc1_weights[113][160] = 16'sd73;
        fc1_weights[113][161] = 16'sd81;
        fc1_weights[113][162] = 16'sd43;
        fc1_weights[113][163] = 16'sd-10;
        fc1_weights[113][164] = 16'sd52;
        fc1_weights[113][165] = 16'sd47;
        fc1_weights[113][166] = 16'sd16;
        fc1_weights[113][167] = 16'sd12;
        fc1_weights[113][168] = 16'sd41;
        fc1_weights[113][169] = 16'sd43;
        fc1_weights[113][170] = 16'sd29;
        fc1_weights[113][171] = 16'sd57;
        fc1_weights[113][172] = 16'sd79;
        fc1_weights[113][173] = 16'sd53;
        fc1_weights[113][174] = 16'sd45;
        fc1_weights[113][175] = 16'sd36;
        fc1_weights[113][176] = 16'sd4;
        fc1_weights[113][177] = 16'sd-96;
        fc1_weights[113][178] = 16'sd2;
        fc1_weights[113][179] = 16'sd30;
        fc1_weights[113][180] = 16'sd-96;
        fc1_weights[113][181] = 16'sd21;
        fc1_weights[113][182] = 16'sd51;
        fc1_weights[113][183] = 16'sd18;
        fc1_weights[113][184] = 16'sd27;
        fc1_weights[113][185] = 16'sd16;
        fc1_weights[113][186] = 16'sd48;
        fc1_weights[113][187] = 16'sd4;
        fc1_weights[113][188] = 16'sd26;
        fc1_weights[113][189] = 16'sd56;
        fc1_weights[113][190] = 16'sd33;
        fc1_weights[113][191] = 16'sd-34;
        fc1_weights[113][192] = 16'sd4;
        fc1_weights[113][193] = 16'sd45;
        fc1_weights[113][194] = 16'sd17;
        fc1_weights[113][195] = 16'sd62;
        fc1_weights[113][196] = 16'sd30;
        fc1_weights[113][197] = 16'sd10;
        fc1_weights[113][198] = 16'sd31;
        fc1_weights[113][199] = 16'sd-37;
        fc1_weights[113][200] = 16'sd2;
        fc1_weights[113][201] = 16'sd30;
        fc1_weights[113][202] = 16'sd-52;
        fc1_weights[113][203] = 16'sd-80;
        fc1_weights[113][204] = 16'sd-34;
        fc1_weights[113][205] = 16'sd-81;
        fc1_weights[113][206] = 16'sd-65;
        fc1_weights[113][207] = 16'sd23;
        fc1_weights[114][0] = 16'sd-57;
        fc1_weights[114][1] = 16'sd19;
        fc1_weights[114][2] = 16'sd-31;
        fc1_weights[114][3] = 16'sd-36;
        fc1_weights[114][4] = 16'sd-18;
        fc1_weights[114][5] = 16'sd23;
        fc1_weights[114][6] = 16'sd-1;
        fc1_weights[114][7] = 16'sd72;
        fc1_weights[114][8] = 16'sd-74;
        fc1_weights[114][9] = 16'sd10;
        fc1_weights[114][10] = 16'sd-11;
        fc1_weights[114][11] = 16'sd-3;
        fc1_weights[114][12] = 16'sd23;
        fc1_weights[114][13] = 16'sd85;
        fc1_weights[114][14] = 16'sd67;
        fc1_weights[114][15] = 16'sd12;
        fc1_weights[114][16] = 16'sd58;
        fc1_weights[114][17] = 16'sd53;
        fc1_weights[114][18] = 16'sd60;
        fc1_weights[114][19] = 16'sd-17;
        fc1_weights[114][20] = 16'sd3;
        fc1_weights[114][21] = 16'sd0;
        fc1_weights[114][22] = 16'sd-7;
        fc1_weights[114][23] = 16'sd18;
        fc1_weights[114][24] = 16'sd-12;
        fc1_weights[114][25] = 16'sd52;
        fc1_weights[114][26] = 16'sd-79;
        fc1_weights[114][27] = 16'sd-47;
        fc1_weights[114][28] = 16'sd-48;
        fc1_weights[114][29] = 16'sd41;
        fc1_weights[114][30] = 16'sd26;
        fc1_weights[114][31] = 16'sd-4;
        fc1_weights[114][32] = 16'sd43;
        fc1_weights[114][33] = 16'sd-57;
        fc1_weights[114][34] = 16'sd25;
        fc1_weights[114][35] = 16'sd-1;
        fc1_weights[114][36] = 16'sd46;
        fc1_weights[114][37] = 16'sd9;
        fc1_weights[114][38] = 16'sd32;
        fc1_weights[114][39] = 16'sd71;
        fc1_weights[114][40] = 16'sd94;
        fc1_weights[114][41] = 16'sd-5;
        fc1_weights[114][42] = 16'sd-24;
        fc1_weights[114][43] = 16'sd-33;
        fc1_weights[114][44] = 16'sd-58;
        fc1_weights[114][45] = 16'sd-22;
        fc1_weights[114][46] = 16'sd-10;
        fc1_weights[114][47] = 16'sd-11;
        fc1_weights[114][48] = 16'sd-34;
        fc1_weights[114][49] = 16'sd10;
        fc1_weights[114][50] = 16'sd-35;
        fc1_weights[114][51] = 16'sd-54;
        fc1_weights[114][52] = 16'sd-17;
        fc1_weights[114][53] = 16'sd-74;
        fc1_weights[114][54] = 16'sd-21;
        fc1_weights[114][55] = 16'sd-3;
        fc1_weights[114][56] = 16'sd39;
        fc1_weights[114][57] = 16'sd-33;
        fc1_weights[114][58] = 16'sd-19;
        fc1_weights[114][59] = 16'sd-56;
        fc1_weights[114][60] = 16'sd49;
        fc1_weights[114][61] = 16'sd42;
        fc1_weights[114][62] = 16'sd-25;
        fc1_weights[114][63] = 16'sd64;
        fc1_weights[114][64] = 16'sd64;
        fc1_weights[114][65] = 16'sd-45;
        fc1_weights[114][66] = 16'sd61;
        fc1_weights[114][67] = 16'sd-10;
        fc1_weights[114][68] = 16'sd-76;
        fc1_weights[114][69] = 16'sd28;
        fc1_weights[114][70] = 16'sd-35;
        fc1_weights[114][71] = 16'sd8;
        fc1_weights[114][72] = 16'sd0;
        fc1_weights[114][73] = 16'sd21;
        fc1_weights[114][74] = 16'sd62;
        fc1_weights[114][75] = 16'sd1;
        fc1_weights[114][76] = 16'sd33;
        fc1_weights[114][77] = 16'sd0;
        fc1_weights[114][78] = 16'sd-17;
        fc1_weights[114][79] = 16'sd6;
        fc1_weights[114][80] = 16'sd-20;
        fc1_weights[114][81] = 16'sd-72;
        fc1_weights[114][82] = 16'sd-51;
        fc1_weights[114][83] = 16'sd-36;
        fc1_weights[114][84] = 16'sd6;
        fc1_weights[114][85] = 16'sd-34;
        fc1_weights[114][86] = 16'sd-24;
        fc1_weights[114][87] = 16'sd19;
        fc1_weights[114][88] = 16'sd-29;
        fc1_weights[114][89] = 16'sd-76;
        fc1_weights[114][90] = 16'sd-20;
        fc1_weights[114][91] = 16'sd50;
        fc1_weights[114][92] = 16'sd33;
        fc1_weights[114][93] = 16'sd-16;
        fc1_weights[114][94] = 16'sd-44;
        fc1_weights[114][95] = 16'sd56;
        fc1_weights[114][96] = 16'sd-7;
        fc1_weights[114][97] = 16'sd-17;
        fc1_weights[114][98] = 16'sd13;
        fc1_weights[114][99] = 16'sd-41;
        fc1_weights[114][100] = 16'sd52;
        fc1_weights[114][101] = 16'sd-15;
        fc1_weights[114][102] = 16'sd-28;
        fc1_weights[114][103] = 16'sd-6;
        fc1_weights[114][104] = 16'sd5;
        fc1_weights[114][105] = 16'sd-87;
        fc1_weights[114][106] = 16'sd35;
        fc1_weights[114][107] = 16'sd-47;
        fc1_weights[114][108] = 16'sd-18;
        fc1_weights[114][109] = 16'sd-19;
        fc1_weights[114][110] = 16'sd12;
        fc1_weights[114][111] = 16'sd-18;
        fc1_weights[114][112] = 16'sd27;
        fc1_weights[114][113] = 16'sd-25;
        fc1_weights[114][114] = 16'sd7;
        fc1_weights[114][115] = 16'sd-14;
        fc1_weights[114][116] = 16'sd9;
        fc1_weights[114][117] = 16'sd31;
        fc1_weights[114][118] = 16'sd29;
        fc1_weights[114][119] = 16'sd15;
        fc1_weights[114][120] = 16'sd-20;
        fc1_weights[114][121] = 16'sd9;
        fc1_weights[114][122] = 16'sd-2;
        fc1_weights[114][123] = 16'sd-12;
        fc1_weights[114][124] = 16'sd17;
        fc1_weights[114][125] = 16'sd-30;
        fc1_weights[114][126] = 16'sd-12;
        fc1_weights[114][127] = 16'sd-12;
        fc1_weights[114][128] = 16'sd46;
        fc1_weights[114][129] = 16'sd59;
        fc1_weights[114][130] = 16'sd2;
        fc1_weights[114][131] = 16'sd45;
        fc1_weights[114][132] = 16'sd28;
        fc1_weights[114][133] = 16'sd-2;
        fc1_weights[114][134] = 16'sd24;
        fc1_weights[114][135] = 16'sd39;
        fc1_weights[114][136] = 16'sd38;
        fc1_weights[114][137] = 16'sd-4;
        fc1_weights[114][138] = 16'sd41;
        fc1_weights[114][139] = 16'sd-20;
        fc1_weights[114][140] = 16'sd20;
        fc1_weights[114][141] = 16'sd10;
        fc1_weights[114][142] = 16'sd22;
        fc1_weights[114][143] = 16'sd-12;
        fc1_weights[114][144] = 16'sd68;
        fc1_weights[114][145] = 16'sd-13;
        fc1_weights[114][146] = 16'sd3;
        fc1_weights[114][147] = 16'sd-5;
        fc1_weights[114][148] = 16'sd-13;
        fc1_weights[114][149] = 16'sd-29;
        fc1_weights[114][150] = 16'sd-22;
        fc1_weights[114][151] = 16'sd-18;
        fc1_weights[114][152] = 16'sd15;
        fc1_weights[114][153] = 16'sd-13;
        fc1_weights[114][154] = 16'sd70;
        fc1_weights[114][155] = 16'sd-10;
        fc1_weights[114][156] = 16'sd9;
        fc1_weights[114][157] = 16'sd0;
        fc1_weights[114][158] = 16'sd6;
        fc1_weights[114][159] = 16'sd15;
        fc1_weights[114][160] = 16'sd-44;
        fc1_weights[114][161] = 16'sd2;
        fc1_weights[114][162] = 16'sd-2;
        fc1_weights[114][163] = 16'sd0;
        fc1_weights[114][164] = 16'sd13;
        fc1_weights[114][165] = 16'sd3;
        fc1_weights[114][166] = 16'sd-64;
        fc1_weights[114][167] = 16'sd-37;
        fc1_weights[114][168] = 16'sd-25;
        fc1_weights[114][169] = 16'sd-27;
        fc1_weights[114][170] = 16'sd16;
        fc1_weights[114][171] = 16'sd-51;
        fc1_weights[114][172] = 16'sd-42;
        fc1_weights[114][173] = 16'sd-54;
        fc1_weights[114][174] = 16'sd-26;
        fc1_weights[114][175] = 16'sd-53;
        fc1_weights[114][176] = 16'sd-63;
        fc1_weights[114][177] = 16'sd18;
        fc1_weights[114][178] = 16'sd13;
        fc1_weights[114][179] = 16'sd-20;
        fc1_weights[114][180] = 16'sd-29;
        fc1_weights[114][181] = 16'sd-15;
        fc1_weights[114][182] = 16'sd36;
        fc1_weights[114][183] = 16'sd18;
        fc1_weights[114][184] = 16'sd48;
        fc1_weights[114][185] = 16'sd19;
        fc1_weights[114][186] = 16'sd-29;
        fc1_weights[114][187] = 16'sd-30;
        fc1_weights[114][188] = 16'sd-32;
        fc1_weights[114][189] = 16'sd-34;
        fc1_weights[114][190] = 16'sd34;
        fc1_weights[114][191] = 16'sd-6;
        fc1_weights[114][192] = 16'sd18;
        fc1_weights[114][193] = 16'sd-25;
        fc1_weights[114][194] = 16'sd22;
        fc1_weights[114][195] = 16'sd0;
        fc1_weights[114][196] = 16'sd-20;
        fc1_weights[114][197] = 16'sd-24;
        fc1_weights[114][198] = 16'sd3;
        fc1_weights[114][199] = 16'sd-70;
        fc1_weights[114][200] = 16'sd16;
        fc1_weights[114][201] = 16'sd-28;
        fc1_weights[114][202] = 16'sd-4;
        fc1_weights[114][203] = 16'sd52;
        fc1_weights[114][204] = 16'sd-13;
        fc1_weights[114][205] = 16'sd-8;
        fc1_weights[114][206] = 16'sd46;
        fc1_weights[114][207] = 16'sd67;
        fc1_weights[115][0] = 16'sd-33;
        fc1_weights[115][1] = 16'sd-30;
        fc1_weights[115][2] = 16'sd-23;
        fc1_weights[115][3] = 16'sd-74;
        fc1_weights[115][4] = 16'sd6;
        fc1_weights[115][5] = 16'sd7;
        fc1_weights[115][6] = 16'sd40;
        fc1_weights[115][7] = 16'sd-5;
        fc1_weights[115][8] = 16'sd-6;
        fc1_weights[115][9] = 16'sd-32;
        fc1_weights[115][10] = 16'sd-93;
        fc1_weights[115][11] = 16'sd-34;
        fc1_weights[115][12] = 16'sd33;
        fc1_weights[115][13] = 16'sd38;
        fc1_weights[115][14] = 16'sd1;
        fc1_weights[115][15] = 16'sd-3;
        fc1_weights[115][16] = 16'sd-3;
        fc1_weights[115][17] = 16'sd59;
        fc1_weights[115][18] = 16'sd44;
        fc1_weights[115][19] = 16'sd11;
        fc1_weights[115][20] = 16'sd32;
        fc1_weights[115][21] = 16'sd-17;
        fc1_weights[115][22] = 16'sd1;
        fc1_weights[115][23] = 16'sd58;
        fc1_weights[115][24] = 16'sd9;
        fc1_weights[115][25] = 16'sd41;
        fc1_weights[115][26] = 16'sd-9;
        fc1_weights[115][27] = 16'sd18;
        fc1_weights[115][28] = 16'sd-20;
        fc1_weights[115][29] = 16'sd-45;
        fc1_weights[115][30] = 16'sd-41;
        fc1_weights[115][31] = 16'sd-42;
        fc1_weights[115][32] = 16'sd20;
        fc1_weights[115][33] = 16'sd38;
        fc1_weights[115][34] = 16'sd32;
        fc1_weights[115][35] = 16'sd-11;
        fc1_weights[115][36] = 16'sd-54;
        fc1_weights[115][37] = 16'sd-47;
        fc1_weights[115][38] = 16'sd-30;
        fc1_weights[115][39] = 16'sd-34;
        fc1_weights[115][40] = 16'sd-68;
        fc1_weights[115][41] = 16'sd52;
        fc1_weights[115][42] = 16'sd-1;
        fc1_weights[115][43] = 16'sd-23;
        fc1_weights[115][44] = 16'sd6;
        fc1_weights[115][45] = 16'sd54;
        fc1_weights[115][46] = 16'sd24;
        fc1_weights[115][47] = 16'sd8;
        fc1_weights[115][48] = 16'sd-11;
        fc1_weights[115][49] = 16'sd11;
        fc1_weights[115][50] = 16'sd22;
        fc1_weights[115][51] = 16'sd77;
        fc1_weights[115][52] = 16'sd-15;
        fc1_weights[115][53] = 16'sd-16;
        fc1_weights[115][54] = 16'sd-51;
        fc1_weights[115][55] = 16'sd-48;
        fc1_weights[115][56] = 16'sd-24;
        fc1_weights[115][57] = 16'sd-59;
        fc1_weights[115][58] = 16'sd1;
        fc1_weights[115][59] = 16'sd3;
        fc1_weights[115][60] = 16'sd-39;
        fc1_weights[115][61] = 16'sd5;
        fc1_weights[115][62] = 16'sd35;
        fc1_weights[115][63] = 16'sd11;
        fc1_weights[115][64] = 16'sd41;
        fc1_weights[115][65] = 16'sd-16;
        fc1_weights[115][66] = 16'sd-28;
        fc1_weights[115][67] = 16'sd-16;
        fc1_weights[115][68] = 16'sd7;
        fc1_weights[115][69] = 16'sd-36;
        fc1_weights[115][70] = 16'sd11;
        fc1_weights[115][71] = 16'sd33;
        fc1_weights[115][72] = 16'sd-15;
        fc1_weights[115][73] = 16'sd42;
        fc1_weights[115][74] = 16'sd11;
        fc1_weights[115][75] = 16'sd-5;
        fc1_weights[115][76] = 16'sd-50;
        fc1_weights[115][77] = 16'sd20;
        fc1_weights[115][78] = 16'sd-14;
        fc1_weights[115][79] = 16'sd-24;
        fc1_weights[115][80] = 16'sd-10;
        fc1_weights[115][81] = 16'sd17;
        fc1_weights[115][82] = 16'sd10;
        fc1_weights[115][83] = 16'sd-7;
        fc1_weights[115][84] = 16'sd-8;
        fc1_weights[115][85] = 16'sd89;
        fc1_weights[115][86] = 16'sd12;
        fc1_weights[115][87] = 16'sd0;
        fc1_weights[115][88] = 16'sd70;
        fc1_weights[115][89] = 16'sd-25;
        fc1_weights[115][90] = 16'sd-2;
        fc1_weights[115][91] = 16'sd-34;
        fc1_weights[115][92] = 16'sd-77;
        fc1_weights[115][93] = 16'sd-45;
        fc1_weights[115][94] = 16'sd-45;
        fc1_weights[115][95] = 16'sd-39;
        fc1_weights[115][96] = 16'sd-28;
        fc1_weights[115][97] = 16'sd-49;
        fc1_weights[115][98] = 16'sd-21;
        fc1_weights[115][99] = 16'sd-40;
        fc1_weights[115][100] = 16'sd-13;
        fc1_weights[115][101] = 16'sd-21;
        fc1_weights[115][102] = 16'sd-13;
        fc1_weights[115][103] = 16'sd-1;
        fc1_weights[115][104] = 16'sd-1;
        fc1_weights[115][105] = 16'sd-24;
        fc1_weights[115][106] = 16'sd-7;
        fc1_weights[115][107] = 16'sd33;
        fc1_weights[115][108] = 16'sd-21;
        fc1_weights[115][109] = 16'sd-1;
        fc1_weights[115][110] = 16'sd-22;
        fc1_weights[115][111] = 16'sd-36;
        fc1_weights[115][112] = 16'sd-3;
        fc1_weights[115][113] = 16'sd0;
        fc1_weights[115][114] = 16'sd-16;
        fc1_weights[115][115] = 16'sd-8;
        fc1_weights[115][116] = 16'sd7;
        fc1_weights[115][117] = 16'sd57;
        fc1_weights[115][118] = 16'sd-13;
        fc1_weights[115][119] = 16'sd17;
        fc1_weights[115][120] = 16'sd24;
        fc1_weights[115][121] = 16'sd-21;
        fc1_weights[115][122] = 16'sd-66;
        fc1_weights[115][123] = 16'sd-14;
        fc1_weights[115][124] = 16'sd-6;
        fc1_weights[115][125] = 16'sd-14;
        fc1_weights[115][126] = 16'sd25;
        fc1_weights[115][127] = 16'sd-31;
        fc1_weights[115][128] = 16'sd-2;
        fc1_weights[115][129] = 16'sd14;
        fc1_weights[115][130] = 16'sd11;
        fc1_weights[115][131] = 16'sd23;
        fc1_weights[115][132] = 16'sd5;
        fc1_weights[115][133] = 16'sd-15;
        fc1_weights[115][134] = 16'sd-17;
        fc1_weights[115][135] = 16'sd-44;
        fc1_weights[115][136] = 16'sd-10;
        fc1_weights[115][137] = 16'sd-20;
        fc1_weights[115][138] = 16'sd-57;
        fc1_weights[115][139] = 16'sd-20;
        fc1_weights[115][140] = 16'sd-39;
        fc1_weights[115][141] = 16'sd-6;
        fc1_weights[115][142] = 16'sd-34;
        fc1_weights[115][143] = 16'sd21;
        fc1_weights[115][144] = 16'sd34;
        fc1_weights[115][145] = 16'sd12;
        fc1_weights[115][146] = 16'sd12;
        fc1_weights[115][147] = 16'sd-2;
        fc1_weights[115][148] = 16'sd-45;
        fc1_weights[115][149] = 16'sd-26;
        fc1_weights[115][150] = 16'sd-28;
        fc1_weights[115][151] = 16'sd-12;
        fc1_weights[115][152] = 16'sd-3;
        fc1_weights[115][153] = 16'sd-20;
        fc1_weights[115][154] = 16'sd-42;
        fc1_weights[115][155] = 16'sd-4;
        fc1_weights[115][156] = 16'sd-18;
        fc1_weights[115][157] = 16'sd-18;
        fc1_weights[115][158] = 16'sd-7;
        fc1_weights[115][159] = 16'sd16;
        fc1_weights[115][160] = 16'sd4;
        fc1_weights[115][161] = 16'sd-33;
        fc1_weights[115][162] = 16'sd-65;
        fc1_weights[115][163] = 16'sd-31;
        fc1_weights[115][164] = 16'sd25;
        fc1_weights[115][165] = 16'sd18;
        fc1_weights[115][166] = 16'sd-29;
        fc1_weights[115][167] = 16'sd-43;
        fc1_weights[115][168] = 16'sd-46;
        fc1_weights[115][169] = 16'sd8;
        fc1_weights[115][170] = 16'sd18;
        fc1_weights[115][171] = 16'sd-29;
        fc1_weights[115][172] = 16'sd-27;
        fc1_weights[115][173] = 16'sd-16;
        fc1_weights[115][174] = 16'sd22;
        fc1_weights[115][175] = 16'sd22;
        fc1_weights[115][176] = 16'sd7;
        fc1_weights[115][177] = 16'sd16;
        fc1_weights[115][178] = 16'sd31;
        fc1_weights[115][179] = 16'sd-26;
        fc1_weights[115][180] = 16'sd37;
        fc1_weights[115][181] = 16'sd14;
        fc1_weights[115][182] = 16'sd-12;
        fc1_weights[115][183] = 16'sd-4;
        fc1_weights[115][184] = 16'sd28;
        fc1_weights[115][185] = 16'sd-30;
        fc1_weights[115][186] = 16'sd-28;
        fc1_weights[115][187] = 16'sd-12;
        fc1_weights[115][188] = 16'sd-3;
        fc1_weights[115][189] = 16'sd37;
        fc1_weights[115][190] = 16'sd51;
        fc1_weights[115][191] = 16'sd-47;
        fc1_weights[115][192] = 16'sd20;
        fc1_weights[115][193] = 16'sd-24;
        fc1_weights[115][194] = 16'sd-8;
        fc1_weights[115][195] = 16'sd1;
        fc1_weights[115][196] = 16'sd44;
        fc1_weights[115][197] = 16'sd-27;
        fc1_weights[115][198] = 16'sd-9;
        fc1_weights[115][199] = 16'sd18;
        fc1_weights[115][200] = 16'sd18;
        fc1_weights[115][201] = 16'sd9;
        fc1_weights[115][202] = 16'sd4;
        fc1_weights[115][203] = 16'sd43;
        fc1_weights[115][204] = 16'sd-26;
        fc1_weights[115][205] = 16'sd39;
        fc1_weights[115][206] = 16'sd78;
        fc1_weights[115][207] = 16'sd88;
        fc1_weights[116][0] = 16'sd9;
        fc1_weights[116][1] = 16'sd-53;
        fc1_weights[116][2] = 16'sd-30;
        fc1_weights[116][3] = 16'sd12;
        fc1_weights[116][4] = 16'sd3;
        fc1_weights[116][5] = 16'sd-13;
        fc1_weights[116][6] = 16'sd17;
        fc1_weights[116][7] = 16'sd-24;
        fc1_weights[116][8] = 16'sd-40;
        fc1_weights[116][9] = 16'sd-41;
        fc1_weights[116][10] = 16'sd0;
        fc1_weights[116][11] = 16'sd-3;
        fc1_weights[116][12] = 16'sd-59;
        fc1_weights[116][13] = 16'sd-69;
        fc1_weights[116][14] = 16'sd-63;
        fc1_weights[116][15] = 16'sd27;
        fc1_weights[116][16] = 16'sd-25;
        fc1_weights[116][17] = 16'sd-19;
        fc1_weights[116][18] = 16'sd-5;
        fc1_weights[116][19] = 16'sd-29;
        fc1_weights[116][20] = 16'sd-13;
        fc1_weights[116][21] = 16'sd-7;
        fc1_weights[116][22] = 16'sd-20;
        fc1_weights[116][23] = 16'sd-45;
        fc1_weights[116][24] = 16'sd-25;
        fc1_weights[116][25] = 16'sd-21;
        fc1_weights[116][26] = 16'sd38;
        fc1_weights[116][27] = 16'sd-24;
        fc1_weights[116][28] = 16'sd-11;
        fc1_weights[116][29] = 16'sd-35;
        fc1_weights[116][30] = 16'sd12;
        fc1_weights[116][31] = 16'sd15;
        fc1_weights[116][32] = 16'sd-10;
        fc1_weights[116][33] = 16'sd-5;
        fc1_weights[116][34] = 16'sd-30;
        fc1_weights[116][35] = 16'sd-50;
        fc1_weights[116][36] = 16'sd-3;
        fc1_weights[116][37] = 16'sd-2;
        fc1_weights[116][38] = 16'sd32;
        fc1_weights[116][39] = 16'sd-69;
        fc1_weights[116][40] = 16'sd20;
        fc1_weights[116][41] = 16'sd17;
        fc1_weights[116][42] = 16'sd-5;
        fc1_weights[116][43] = 16'sd43;
        fc1_weights[116][44] = 16'sd33;
        fc1_weights[116][45] = 16'sd-4;
        fc1_weights[116][46] = 16'sd50;
        fc1_weights[116][47] = 16'sd-18;
        fc1_weights[116][48] = 16'sd47;
        fc1_weights[116][49] = 16'sd43;
        fc1_weights[116][50] = 16'sd4;
        fc1_weights[116][51] = 16'sd16;
        fc1_weights[116][52] = 16'sd0;
        fc1_weights[116][53] = 16'sd41;
        fc1_weights[116][54] = 16'sd-13;
        fc1_weights[116][55] = 16'sd-26;
        fc1_weights[116][56] = 16'sd-41;
        fc1_weights[116][57] = 16'sd-20;
        fc1_weights[116][58] = 16'sd-58;
        fc1_weights[116][59] = 16'sd-29;
        fc1_weights[116][60] = 16'sd-9;
        fc1_weights[116][61] = 16'sd-52;
        fc1_weights[116][62] = 16'sd-18;
        fc1_weights[116][63] = 16'sd0;
        fc1_weights[116][64] = 16'sd-42;
        fc1_weights[116][65] = 16'sd35;
        fc1_weights[116][66] = 16'sd40;
        fc1_weights[116][67] = 16'sd51;
        fc1_weights[116][68] = 16'sd20;
        fc1_weights[116][69] = 16'sd27;
        fc1_weights[116][70] = 16'sd-26;
        fc1_weights[116][71] = 16'sd-38;
        fc1_weights[116][72] = 16'sd-21;
        fc1_weights[116][73] = 16'sd-28;
        fc1_weights[116][74] = 16'sd-11;
        fc1_weights[116][75] = 16'sd22;
        fc1_weights[116][76] = 16'sd54;
        fc1_weights[116][77] = 16'sd20;
        fc1_weights[116][78] = 16'sd38;
        fc1_weights[116][79] = 16'sd55;
        fc1_weights[116][80] = 16'sd17;
        fc1_weights[116][81] = 16'sd22;
        fc1_weights[116][82] = 16'sd27;
        fc1_weights[116][83] = 16'sd-65;
        fc1_weights[116][84] = 16'sd-23;
        fc1_weights[116][85] = 16'sd-23;
        fc1_weights[116][86] = 16'sd-30;
        fc1_weights[116][87] = 16'sd-73;
        fc1_weights[116][88] = 16'sd-48;
        fc1_weights[116][89] = 16'sd61;
        fc1_weights[116][90] = 16'sd5;
        fc1_weights[116][91] = 16'sd39;
        fc1_weights[116][92] = 16'sd49;
        fc1_weights[116][93] = 16'sd118;
        fc1_weights[116][94] = 16'sd69;
        fc1_weights[116][95] = 16'sd-6;
        fc1_weights[116][96] = 16'sd-2;
        fc1_weights[116][97] = 16'sd20;
        fc1_weights[116][98] = 16'sd-6;
        fc1_weights[116][99] = 16'sd32;
        fc1_weights[116][100] = 16'sd14;
        fc1_weights[116][101] = 16'sd71;
        fc1_weights[116][102] = 16'sd43;
        fc1_weights[116][103] = 16'sd5;
        fc1_weights[116][104] = 16'sd-8;
        fc1_weights[116][105] = 16'sd25;
        fc1_weights[116][106] = 16'sd-7;
        fc1_weights[116][107] = 16'sd24;
        fc1_weights[116][108] = 16'sd12;
        fc1_weights[116][109] = 16'sd5;
        fc1_weights[116][110] = 16'sd-9;
        fc1_weights[116][111] = 16'sd-33;
        fc1_weights[116][112] = 16'sd32;
        fc1_weights[116][113] = 16'sd-12;
        fc1_weights[116][114] = 16'sd10;
        fc1_weights[116][115] = 16'sd-9;
        fc1_weights[116][116] = 16'sd41;
        fc1_weights[116][117] = 16'sd57;
        fc1_weights[116][118] = 16'sd1;
        fc1_weights[116][119] = 16'sd65;
        fc1_weights[116][120] = 16'sd15;
        fc1_weights[116][121] = 16'sd20;
        fc1_weights[116][122] = 16'sd-4;
        fc1_weights[116][123] = 16'sd14;
        fc1_weights[116][124] = 16'sd23;
        fc1_weights[116][125] = 16'sd-24;
        fc1_weights[116][126] = 16'sd-43;
        fc1_weights[116][127] = 16'sd0;
        fc1_weights[116][128] = 16'sd14;
        fc1_weights[116][129] = 16'sd-15;
        fc1_weights[116][130] = 16'sd-18;
        fc1_weights[116][131] = 16'sd-30;
        fc1_weights[116][132] = 16'sd-21;
        fc1_weights[116][133] = 16'sd-2;
        fc1_weights[116][134] = 16'sd24;
        fc1_weights[116][135] = 16'sd30;
        fc1_weights[116][136] = 16'sd2;
        fc1_weights[116][137] = 16'sd33;
        fc1_weights[116][138] = 16'sd31;
        fc1_weights[116][139] = 16'sd60;
        fc1_weights[116][140] = 16'sd-28;
        fc1_weights[116][141] = 16'sd-42;
        fc1_weights[116][142] = 16'sd-3;
        fc1_weights[116][143] = 16'sd-50;
        fc1_weights[116][144] = 16'sd25;
        fc1_weights[116][145] = 16'sd4;
        fc1_weights[116][146] = 16'sd39;
        fc1_weights[116][147] = 16'sd22;
        fc1_weights[116][148] = 16'sd40;
        fc1_weights[116][149] = 16'sd41;
        fc1_weights[116][150] = 16'sd16;
        fc1_weights[116][151] = 16'sd-21;
        fc1_weights[116][152] = 16'sd23;
        fc1_weights[116][153] = 16'sd1;
        fc1_weights[116][154] = 16'sd13;
        fc1_weights[116][155] = 16'sd-24;
        fc1_weights[116][156] = 16'sd-12;
        fc1_weights[116][157] = 16'sd-4;
        fc1_weights[116][158] = 16'sd16;
        fc1_weights[116][159] = 16'sd23;
        fc1_weights[116][160] = 16'sd21;
        fc1_weights[116][161] = 16'sd2;
        fc1_weights[116][162] = 16'sd32;
        fc1_weights[116][163] = 16'sd34;
        fc1_weights[116][164] = 16'sd51;
        fc1_weights[116][165] = 16'sd19;
        fc1_weights[116][166] = 16'sd28;
        fc1_weights[116][167] = 16'sd8;
        fc1_weights[116][168] = 16'sd39;
        fc1_weights[116][169] = 16'sd-36;
        fc1_weights[116][170] = 16'sd-38;
        fc1_weights[116][171] = 16'sd-8;
        fc1_weights[116][172] = 16'sd2;
        fc1_weights[116][173] = 16'sd9;
        fc1_weights[116][174] = 16'sd13;
        fc1_weights[116][175] = 16'sd11;
        fc1_weights[116][176] = 16'sd15;
        fc1_weights[116][177] = 16'sd36;
        fc1_weights[116][178] = 16'sd-26;
        fc1_weights[116][179] = 16'sd-9;
        fc1_weights[116][180] = 16'sd22;
        fc1_weights[116][181] = 16'sd13;
        fc1_weights[116][182] = 16'sd-38;
        fc1_weights[116][183] = 16'sd57;
        fc1_weights[116][184] = 16'sd9;
        fc1_weights[116][185] = 16'sd48;
        fc1_weights[116][186] = 16'sd47;
        fc1_weights[116][187] = 16'sd80;
        fc1_weights[116][188] = 16'sd89;
        fc1_weights[116][189] = 16'sd77;
        fc1_weights[116][190] = 16'sd52;
        fc1_weights[116][191] = 16'sd45;
        fc1_weights[116][192] = 16'sd-25;
        fc1_weights[116][193] = 16'sd8;
        fc1_weights[116][194] = 16'sd-2;
        fc1_weights[116][195] = 16'sd3;
        fc1_weights[116][196] = 16'sd-5;
        fc1_weights[116][197] = 16'sd75;
        fc1_weights[116][198] = 16'sd1;
        fc1_weights[116][199] = 16'sd32;
        fc1_weights[116][200] = 16'sd0;
        fc1_weights[116][201] = 16'sd27;
        fc1_weights[116][202] = 16'sd-1;
        fc1_weights[116][203] = 16'sd-17;
        fc1_weights[116][204] = 16'sd30;
        fc1_weights[116][205] = 16'sd72;
        fc1_weights[116][206] = 16'sd-17;
        fc1_weights[116][207] = 16'sd-31;
        fc1_weights[117][0] = 16'sd40;
        fc1_weights[117][1] = 16'sd30;
        fc1_weights[117][2] = 16'sd-13;
        fc1_weights[117][3] = 16'sd26;
        fc1_weights[117][4] = 16'sd-9;
        fc1_weights[117][5] = 16'sd9;
        fc1_weights[117][6] = 16'sd-21;
        fc1_weights[117][7] = 16'sd-17;
        fc1_weights[117][8] = 16'sd20;
        fc1_weights[117][9] = 16'sd62;
        fc1_weights[117][10] = 16'sd4;
        fc1_weights[117][11] = 16'sd20;
        fc1_weights[117][12] = 16'sd-11;
        fc1_weights[117][13] = 16'sd-27;
        fc1_weights[117][14] = 16'sd-54;
        fc1_weights[117][15] = 16'sd-39;
        fc1_weights[117][16] = 16'sd-13;
        fc1_weights[117][17] = 16'sd-13;
        fc1_weights[117][18] = 16'sd-37;
        fc1_weights[117][19] = 16'sd-33;
        fc1_weights[117][20] = 16'sd3;
        fc1_weights[117][21] = 16'sd-23;
        fc1_weights[117][22] = 16'sd4;
        fc1_weights[117][23] = 16'sd17;
        fc1_weights[117][24] = 16'sd-33;
        fc1_weights[117][25] = 16'sd-39;
        fc1_weights[117][26] = 16'sd39;
        fc1_weights[117][27] = 16'sd8;
        fc1_weights[117][28] = 16'sd27;
        fc1_weights[117][29] = 16'sd-46;
        fc1_weights[117][30] = 16'sd-5;
        fc1_weights[117][31] = 16'sd-8;
        fc1_weights[117][32] = 16'sd-11;
        fc1_weights[117][33] = 16'sd42;
        fc1_weights[117][34] = 16'sd-29;
        fc1_weights[117][35] = 16'sd-37;
        fc1_weights[117][36] = 16'sd0;
        fc1_weights[117][37] = 16'sd3;
        fc1_weights[117][38] = 16'sd22;
        fc1_weights[117][39] = 16'sd-55;
        fc1_weights[117][40] = 16'sd-47;
        fc1_weights[117][41] = 16'sd-20;
        fc1_weights[117][42] = 16'sd7;
        fc1_weights[117][43] = 16'sd4;
        fc1_weights[117][44] = 16'sd10;
        fc1_weights[117][45] = 16'sd-24;
        fc1_weights[117][46] = 16'sd-32;
        fc1_weights[117][47] = 16'sd-5;
        fc1_weights[117][48] = 16'sd-13;
        fc1_weights[117][49] = 16'sd-10;
        fc1_weights[117][50] = 16'sd-41;
        fc1_weights[117][51] = 16'sd-45;
        fc1_weights[117][52] = 16'sd14;
        fc1_weights[117][53] = 16'sd-1;
        fc1_weights[117][54] = 16'sd8;
        fc1_weights[117][55] = 16'sd-24;
        fc1_weights[117][56] = 16'sd-25;
        fc1_weights[117][57] = 16'sd-11;
        fc1_weights[117][58] = 16'sd-62;
        fc1_weights[117][59] = 16'sd-35;
        fc1_weights[117][60] = 16'sd-67;
        fc1_weights[117][61] = 16'sd-57;
        fc1_weights[117][62] = 16'sd-46;
        fc1_weights[117][63] = 16'sd0;
        fc1_weights[117][64] = 16'sd-46;
        fc1_weights[117][65] = 16'sd-13;
        fc1_weights[117][66] = 16'sd39;
        fc1_weights[117][67] = 16'sd24;
        fc1_weights[117][68] = 16'sd36;
        fc1_weights[117][69] = 16'sd1;
        fc1_weights[117][70] = 16'sd-74;
        fc1_weights[117][71] = 16'sd20;
        fc1_weights[117][72] = 16'sd14;
        fc1_weights[117][73] = 16'sd-32;
        fc1_weights[117][74] = 16'sd1;
        fc1_weights[117][75] = 16'sd71;
        fc1_weights[117][76] = 16'sd41;
        fc1_weights[117][77] = 16'sd-58;
        fc1_weights[117][78] = 16'sd3;
        fc1_weights[117][79] = 16'sd14;
        fc1_weights[117][80] = 16'sd40;
        fc1_weights[117][81] = 16'sd42;
        fc1_weights[117][82] = 16'sd32;
        fc1_weights[117][83] = 16'sd13;
        fc1_weights[117][84] = 16'sd12;
        fc1_weights[117][85] = 16'sd5;
        fc1_weights[117][86] = 16'sd-10;
        fc1_weights[117][87] = 16'sd-46;
        fc1_weights[117][88] = 16'sd-93;
        fc1_weights[117][89] = 16'sd79;
        fc1_weights[117][90] = 16'sd60;
        fc1_weights[117][91] = 16'sd22;
        fc1_weights[117][92] = 16'sd18;
        fc1_weights[117][93] = 16'sd24;
        fc1_weights[117][94] = 16'sd95;
        fc1_weights[117][95] = 16'sd24;
        fc1_weights[117][96] = 16'sd10;
        fc1_weights[117][97] = 16'sd-10;
        fc1_weights[117][98] = 16'sd34;
        fc1_weights[117][99] = 16'sd63;
        fc1_weights[117][100] = 16'sd56;
        fc1_weights[117][101] = 16'sd4;
        fc1_weights[117][102] = 16'sd72;
        fc1_weights[117][103] = 16'sd28;
        fc1_weights[117][104] = 16'sd-3;
        fc1_weights[117][105] = 16'sd48;
        fc1_weights[117][106] = 16'sd30;
        fc1_weights[117][107] = 16'sd8;
        fc1_weights[117][108] = 16'sd25;
        fc1_weights[117][109] = 16'sd33;
        fc1_weights[117][110] = 16'sd22;
        fc1_weights[117][111] = 16'sd3;
        fc1_weights[117][112] = 16'sd26;
        fc1_weights[117][113] = 16'sd19;
        fc1_weights[117][114] = 16'sd-29;
        fc1_weights[117][115] = 16'sd-49;
        fc1_weights[117][116] = 16'sd26;
        fc1_weights[117][117] = 16'sd36;
        fc1_weights[117][118] = 16'sd28;
        fc1_weights[117][119] = 16'sd85;
        fc1_weights[117][120] = 16'sd108;
        fc1_weights[117][121] = 16'sd73;
        fc1_weights[117][122] = 16'sd89;
        fc1_weights[117][123] = 16'sd-1;
        fc1_weights[117][124] = 16'sd103;
        fc1_weights[117][125] = 16'sd8;
        fc1_weights[117][126] = 16'sd9;
        fc1_weights[117][127] = 16'sd-33;
        fc1_weights[117][128] = 16'sd11;
        fc1_weights[117][129] = 16'sd-23;
        fc1_weights[117][130] = 16'sd4;
        fc1_weights[117][131] = 16'sd8;
        fc1_weights[117][132] = 16'sd62;
        fc1_weights[117][133] = 16'sd36;
        fc1_weights[117][134] = 16'sd-19;
        fc1_weights[117][135] = 16'sd25;
        fc1_weights[117][136] = 16'sd-25;
        fc1_weights[117][137] = 16'sd-6;
        fc1_weights[117][138] = 16'sd-144;
        fc1_weights[117][139] = 16'sd-16;
        fc1_weights[117][140] = 16'sd-26;
        fc1_weights[117][141] = 16'sd-85;
        fc1_weights[117][142] = 16'sd21;
        fc1_weights[117][143] = 16'sd-7;
        fc1_weights[117][144] = 16'sd-54;
        fc1_weights[117][145] = 16'sd-38;
        fc1_weights[117][146] = 16'sd32;
        fc1_weights[117][147] = 16'sd-5;
        fc1_weights[117][148] = 16'sd36;
        fc1_weights[117][149] = 16'sd42;
        fc1_weights[117][150] = 16'sd20;
        fc1_weights[117][151] = 16'sd-76;
        fc1_weights[117][152] = 16'sd0;
        fc1_weights[117][153] = 16'sd-24;
        fc1_weights[117][154] = 16'sd30;
        fc1_weights[117][155] = 16'sd-41;
        fc1_weights[117][156] = 16'sd32;
        fc1_weights[117][157] = 16'sd-14;
        fc1_weights[117][158] = 16'sd0;
        fc1_weights[117][159] = 16'sd-50;
        fc1_weights[117][160] = 16'sd1;
        fc1_weights[117][161] = 16'sd-41;
        fc1_weights[117][162] = 16'sd-63;
        fc1_weights[117][163] = 16'sd-33;
        fc1_weights[117][164] = 16'sd24;
        fc1_weights[117][165] = 16'sd58;
        fc1_weights[117][166] = 16'sd28;
        fc1_weights[117][167] = 16'sd53;
        fc1_weights[117][168] = 16'sd51;
        fc1_weights[117][169] = 16'sd17;
        fc1_weights[117][170] = 16'sd20;
        fc1_weights[117][171] = 16'sd48;
        fc1_weights[117][172] = 16'sd-13;
        fc1_weights[117][173] = 16'sd79;
        fc1_weights[117][174] = 16'sd40;
        fc1_weights[117][175] = 16'sd58;
        fc1_weights[117][176] = 16'sd71;
        fc1_weights[117][177] = 16'sd23;
        fc1_weights[117][178] = 16'sd9;
        fc1_weights[117][179] = 16'sd11;
        fc1_weights[117][180] = 16'sd10;
        fc1_weights[117][181] = 16'sd-18;
        fc1_weights[117][182] = 16'sd-61;
        fc1_weights[117][183] = 16'sd25;
        fc1_weights[117][184] = 16'sd-22;
        fc1_weights[117][185] = 16'sd-15;
        fc1_weights[117][186] = 16'sd-26;
        fc1_weights[117][187] = 16'sd19;
        fc1_weights[117][188] = 16'sd3;
        fc1_weights[117][189] = 16'sd0;
        fc1_weights[117][190] = 16'sd-18;
        fc1_weights[117][191] = 16'sd-8;
        fc1_weights[117][192] = 16'sd-12;
        fc1_weights[117][193] = 16'sd7;
        fc1_weights[117][194] = 16'sd39;
        fc1_weights[117][195] = 16'sd25;
        fc1_weights[117][196] = 16'sd52;
        fc1_weights[117][197] = 16'sd54;
        fc1_weights[117][198] = 16'sd80;
        fc1_weights[117][199] = 16'sd79;
        fc1_weights[117][200] = 16'sd-3;
        fc1_weights[117][201] = 16'sd66;
        fc1_weights[117][202] = 16'sd20;
        fc1_weights[117][203] = 16'sd-32;
        fc1_weights[117][204] = 16'sd36;
        fc1_weights[117][205] = 16'sd5;
        fc1_weights[117][206] = 16'sd-31;
        fc1_weights[117][207] = 16'sd-15;
        fc1_weights[118][0] = 16'sd-24;
        fc1_weights[118][1] = 16'sd20;
        fc1_weights[118][2] = 16'sd26;
        fc1_weights[118][3] = 16'sd-15;
        fc1_weights[118][4] = 16'sd-18;
        fc1_weights[118][5] = 16'sd-19;
        fc1_weights[118][6] = 16'sd24;
        fc1_weights[118][7] = 16'sd49;
        fc1_weights[118][8] = 16'sd30;
        fc1_weights[118][9] = 16'sd15;
        fc1_weights[118][10] = 16'sd51;
        fc1_weights[118][11] = 16'sd-8;
        fc1_weights[118][12] = 16'sd67;
        fc1_weights[118][13] = 16'sd32;
        fc1_weights[118][14] = 16'sd-34;
        fc1_weights[118][15] = 16'sd-41;
        fc1_weights[118][16] = 16'sd-57;
        fc1_weights[118][17] = 16'sd22;
        fc1_weights[118][18] = 16'sd17;
        fc1_weights[118][19] = 16'sd5;
        fc1_weights[118][20] = 16'sd14;
        fc1_weights[118][21] = 16'sd73;
        fc1_weights[118][22] = 16'sd85;
        fc1_weights[118][23] = 16'sd28;
        fc1_weights[118][24] = 16'sd-1;
        fc1_weights[118][25] = 16'sd18;
        fc1_weights[118][26] = 16'sd-23;
        fc1_weights[118][27] = 16'sd-9;
        fc1_weights[118][28] = 16'sd41;
        fc1_weights[118][29] = 16'sd0;
        fc1_weights[118][30] = 16'sd9;
        fc1_weights[118][31] = 16'sd-19;
        fc1_weights[118][32] = 16'sd4;
        fc1_weights[118][33] = 16'sd40;
        fc1_weights[118][34] = 16'sd24;
        fc1_weights[118][35] = 16'sd37;
        fc1_weights[118][36] = 16'sd-19;
        fc1_weights[118][37] = 16'sd79;
        fc1_weights[118][38] = 16'sd20;
        fc1_weights[118][39] = 16'sd-36;
        fc1_weights[118][40] = 16'sd31;
        fc1_weights[118][41] = 16'sd30;
        fc1_weights[118][42] = 16'sd39;
        fc1_weights[118][43] = 16'sd-31;
        fc1_weights[118][44] = 16'sd-18;
        fc1_weights[118][45] = 16'sd-1;
        fc1_weights[118][46] = 16'sd-39;
        fc1_weights[118][47] = 16'sd26;
        fc1_weights[118][48] = 16'sd-47;
        fc1_weights[118][49] = 16'sd-10;
        fc1_weights[118][50] = 16'sd-12;
        fc1_weights[118][51] = 16'sd-52;
        fc1_weights[118][52] = 16'sd62;
        fc1_weights[118][53] = 16'sd-51;
        fc1_weights[118][54] = 16'sd20;
        fc1_weights[118][55] = 16'sd-27;
        fc1_weights[118][56] = 16'sd37;
        fc1_weights[118][57] = 16'sd-5;
        fc1_weights[118][58] = 16'sd30;
        fc1_weights[118][59] = 16'sd52;
        fc1_weights[118][60] = 16'sd25;
        fc1_weights[118][61] = 16'sd-18;
        fc1_weights[118][62] = 16'sd20;
        fc1_weights[118][63] = 16'sd66;
        fc1_weights[118][64] = 16'sd-52;
        fc1_weights[118][65] = 16'sd-2;
        fc1_weights[118][66] = 16'sd55;
        fc1_weights[118][67] = 16'sd-25;
        fc1_weights[118][68] = 16'sd-32;
        fc1_weights[118][69] = 16'sd23;
        fc1_weights[118][70] = 16'sd-9;
        fc1_weights[118][71] = 16'sd42;
        fc1_weights[118][72] = 16'sd0;
        fc1_weights[118][73] = 16'sd29;
        fc1_weights[118][74] = 16'sd40;
        fc1_weights[118][75] = 16'sd37;
        fc1_weights[118][76] = 16'sd-48;
        fc1_weights[118][77] = 16'sd-29;
        fc1_weights[118][78] = 16'sd-12;
        fc1_weights[118][79] = 16'sd9;
        fc1_weights[118][80] = 16'sd-44;
        fc1_weights[118][81] = 16'sd-60;
        fc1_weights[118][82] = 16'sd-11;
        fc1_weights[118][83] = 16'sd54;
        fc1_weights[118][84] = 16'sd61;
        fc1_weights[118][85] = 16'sd0;
        fc1_weights[118][86] = 16'sd36;
        fc1_weights[118][87] = 16'sd-18;
        fc1_weights[118][88] = 16'sd30;
        fc1_weights[118][89] = 16'sd8;
        fc1_weights[118][90] = 16'sd-45;
        fc1_weights[118][91] = 16'sd21;
        fc1_weights[118][92] = 16'sd30;
        fc1_weights[118][93] = 16'sd1;
        fc1_weights[118][94] = 16'sd-10;
        fc1_weights[118][95] = 16'sd9;
        fc1_weights[118][96] = 16'sd-25;
        fc1_weights[118][97] = 16'sd-44;
        fc1_weights[118][98] = 16'sd-34;
        fc1_weights[118][99] = 16'sd-46;
        fc1_weights[118][100] = 16'sd5;
        fc1_weights[118][101] = 16'sd-1;
        fc1_weights[118][102] = 16'sd-58;
        fc1_weights[118][103] = 16'sd-28;
        fc1_weights[118][104] = 16'sd102;
        fc1_weights[118][105] = 16'sd22;
        fc1_weights[118][106] = 16'sd20;
        fc1_weights[118][107] = 16'sd-1;
        fc1_weights[118][108] = 16'sd-41;
        fc1_weights[118][109] = 16'sd-49;
        fc1_weights[118][110] = 16'sd-50;
        fc1_weights[118][111] = 16'sd0;
        fc1_weights[118][112] = 16'sd1;
        fc1_weights[118][113] = 16'sd-59;
        fc1_weights[118][114] = 16'sd44;
        fc1_weights[118][115] = 16'sd108;
        fc1_weights[118][116] = 16'sd32;
        fc1_weights[118][117] = 16'sd-17;
        fc1_weights[118][118] = 16'sd-34;
        fc1_weights[118][119] = 16'sd-34;
        fc1_weights[118][120] = 16'sd-2;
        fc1_weights[118][121] = 16'sd-19;
        fc1_weights[118][122] = 16'sd-1;
        fc1_weights[118][123] = 16'sd-82;
        fc1_weights[118][124] = 16'sd-37;
        fc1_weights[118][125] = 16'sd-66;
        fc1_weights[118][126] = 16'sd-12;
        fc1_weights[118][127] = 16'sd-31;
        fc1_weights[118][128] = 16'sd-17;
        fc1_weights[118][129] = 16'sd20;
        fc1_weights[118][130] = 16'sd3;
        fc1_weights[118][131] = 16'sd-6;
        fc1_weights[118][132] = 16'sd-23;
        fc1_weights[118][133] = 16'sd-54;
        fc1_weights[118][134] = 16'sd-38;
        fc1_weights[118][135] = 16'sd-10;
        fc1_weights[118][136] = 16'sd-17;
        fc1_weights[118][137] = 16'sd23;
        fc1_weights[118][138] = 16'sd11;
        fc1_weights[118][139] = 16'sd-33;
        fc1_weights[118][140] = 16'sd60;
        fc1_weights[118][141] = 16'sd141;
        fc1_weights[118][142] = 16'sd-43;
        fc1_weights[118][143] = 16'sd-13;
        fc1_weights[118][144] = 16'sd19;
        fc1_weights[118][145] = 16'sd75;
        fc1_weights[118][146] = 16'sd22;
        fc1_weights[118][147] = 16'sd-31;
        fc1_weights[118][148] = 16'sd-32;
        fc1_weights[118][149] = 16'sd-31;
        fc1_weights[118][150] = 16'sd-25;
        fc1_weights[118][151] = 16'sd-70;
        fc1_weights[118][152] = 16'sd-30;
        fc1_weights[118][153] = 16'sd-7;
        fc1_weights[118][154] = 16'sd51;
        fc1_weights[118][155] = 16'sd-88;
        fc1_weights[118][156] = 16'sd-15;
        fc1_weights[118][157] = 16'sd-30;
        fc1_weights[118][158] = 16'sd77;
        fc1_weights[118][159] = 16'sd95;
        fc1_weights[118][160] = 16'sd35;
        fc1_weights[118][161] = 16'sd31;
        fc1_weights[118][162] = 16'sd31;
        fc1_weights[118][163] = 16'sd-48;
        fc1_weights[118][164] = 16'sd15;
        fc1_weights[118][165] = 16'sd0;
        fc1_weights[118][166] = 16'sd32;
        fc1_weights[118][167] = 16'sd11;
        fc1_weights[118][168] = 16'sd15;
        fc1_weights[118][169] = 16'sd-23;
        fc1_weights[118][170] = 16'sd-88;
        fc1_weights[118][171] = 16'sd-8;
        fc1_weights[118][172] = 16'sd24;
        fc1_weights[118][173] = 16'sd0;
        fc1_weights[118][174] = 16'sd17;
        fc1_weights[118][175] = 16'sd-52;
        fc1_weights[118][176] = 16'sd-46;
        fc1_weights[118][177] = 16'sd-62;
        fc1_weights[118][178] = 16'sd-16;
        fc1_weights[118][179] = 16'sd-44;
        fc1_weights[118][180] = 16'sd-51;
        fc1_weights[118][181] = 16'sd10;
        fc1_weights[118][182] = 16'sd24;
        fc1_weights[118][183] = 16'sd20;
        fc1_weights[118][184] = 16'sd-35;
        fc1_weights[118][185] = 16'sd-24;
        fc1_weights[118][186] = 16'sd-44;
        fc1_weights[118][187] = 16'sd-82;
        fc1_weights[118][188] = 16'sd-11;
        fc1_weights[118][189] = 16'sd-68;
        fc1_weights[118][190] = 16'sd15;
        fc1_weights[118][191] = 16'sd48;
        fc1_weights[118][192] = 16'sd94;
        fc1_weights[118][193] = 16'sd62;
        fc1_weights[118][194] = 16'sd13;
        fc1_weights[118][195] = 16'sd46;
        fc1_weights[118][196] = 16'sd-11;
        fc1_weights[118][197] = 16'sd-73;
        fc1_weights[118][198] = 16'sd13;
        fc1_weights[118][199] = 16'sd69;
        fc1_weights[118][200] = 16'sd41;
        fc1_weights[118][201] = 16'sd39;
        fc1_weights[118][202] = 16'sd-28;
        fc1_weights[118][203] = 16'sd-29;
        fc1_weights[118][204] = 16'sd-50;
        fc1_weights[118][205] = 16'sd-48;
        fc1_weights[118][206] = 16'sd-32;
        fc1_weights[118][207] = 16'sd-17;
        fc1_weights[119][0] = 16'sd-45;
        fc1_weights[119][1] = 16'sd-59;
        fc1_weights[119][2] = 16'sd-19;
        fc1_weights[119][3] = 16'sd-17;
        fc1_weights[119][4] = 16'sd12;
        fc1_weights[119][5] = 16'sd-22;
        fc1_weights[119][6] = 16'sd-13;
        fc1_weights[119][7] = 16'sd8;
        fc1_weights[119][8] = 16'sd22;
        fc1_weights[119][9] = 16'sd25;
        fc1_weights[119][10] = 16'sd-38;
        fc1_weights[119][11] = 16'sd2;
        fc1_weights[119][12] = 16'sd7;
        fc1_weights[119][13] = 16'sd-18;
        fc1_weights[119][14] = 16'sd6;
        fc1_weights[119][15] = 16'sd7;
        fc1_weights[119][16] = 16'sd8;
        fc1_weights[119][17] = 16'sd5;
        fc1_weights[119][18] = 16'sd30;
        fc1_weights[119][19] = 16'sd36;
        fc1_weights[119][20] = 16'sd17;
        fc1_weights[119][21] = 16'sd36;
        fc1_weights[119][22] = 16'sd2;
        fc1_weights[119][23] = 16'sd39;
        fc1_weights[119][24] = 16'sd7;
        fc1_weights[119][25] = 16'sd-9;
        fc1_weights[119][26] = 16'sd-2;
        fc1_weights[119][27] = 16'sd-18;
        fc1_weights[119][28] = 16'sd-7;
        fc1_weights[119][29] = 16'sd-31;
        fc1_weights[119][30] = 16'sd-32;
        fc1_weights[119][31] = 16'sd-54;
        fc1_weights[119][32] = 16'sd-22;
        fc1_weights[119][33] = 16'sd62;
        fc1_weights[119][34] = 16'sd36;
        fc1_weights[119][35] = 16'sd11;
        fc1_weights[119][36] = 16'sd-12;
        fc1_weights[119][37] = 16'sd35;
        fc1_weights[119][38] = 16'sd-10;
        fc1_weights[119][39] = 16'sd17;
        fc1_weights[119][40] = 16'sd-16;
        fc1_weights[119][41] = 16'sd26;
        fc1_weights[119][42] = 16'sd70;
        fc1_weights[119][43] = 16'sd57;
        fc1_weights[119][44] = 16'sd3;
        fc1_weights[119][45] = 16'sd29;
        fc1_weights[119][46] = 16'sd42;
        fc1_weights[119][47] = 16'sd24;
        fc1_weights[119][48] = 16'sd19;
        fc1_weights[119][49] = 16'sd-24;
        fc1_weights[119][50] = 16'sd-2;
        fc1_weights[119][51] = 16'sd38;
        fc1_weights[119][52] = 16'sd-5;
        fc1_weights[119][53] = 16'sd-21;
        fc1_weights[119][54] = 16'sd5;
        fc1_weights[119][55] = 16'sd-14;
        fc1_weights[119][56] = 16'sd26;
        fc1_weights[119][57] = 16'sd8;
        fc1_weights[119][58] = 16'sd5;
        fc1_weights[119][59] = 16'sd14;
        fc1_weights[119][60] = 16'sd-55;
        fc1_weights[119][61] = 16'sd-26;
        fc1_weights[119][62] = 16'sd36;
        fc1_weights[119][63] = 16'sd-25;
        fc1_weights[119][64] = 16'sd-17;
        fc1_weights[119][65] = 16'sd-14;
        fc1_weights[119][66] = 16'sd-21;
        fc1_weights[119][67] = 16'sd56;
        fc1_weights[119][68] = 16'sd42;
        fc1_weights[119][69] = 16'sd5;
        fc1_weights[119][70] = 16'sd12;
        fc1_weights[119][71] = 16'sd49;
        fc1_weights[119][72] = 16'sd11;
        fc1_weights[119][73] = 16'sd7;
        fc1_weights[119][74] = 16'sd6;
        fc1_weights[119][75] = 16'sd-17;
        fc1_weights[119][76] = 16'sd-28;
        fc1_weights[119][77] = 16'sd21;
        fc1_weights[119][78] = 16'sd-1;
        fc1_weights[119][79] = 16'sd-30;
        fc1_weights[119][80] = 16'sd-19;
        fc1_weights[119][81] = 16'sd28;
        fc1_weights[119][82] = 16'sd-23;
        fc1_weights[119][83] = 16'sd21;
        fc1_weights[119][84] = 16'sd53;
        fc1_weights[119][85] = 16'sd56;
        fc1_weights[119][86] = 16'sd7;
        fc1_weights[119][87] = 16'sd2;
        fc1_weights[119][88] = 16'sd28;
        fc1_weights[119][89] = 16'sd26;
        fc1_weights[119][90] = 16'sd-49;
        fc1_weights[119][91] = 16'sd-35;
        fc1_weights[119][92] = 16'sd-50;
        fc1_weights[119][93] = 16'sd-32;
        fc1_weights[119][94] = 16'sd-12;
        fc1_weights[119][95] = 16'sd-41;
        fc1_weights[119][96] = 16'sd-19;
        fc1_weights[119][97] = 16'sd21;
        fc1_weights[119][98] = 16'sd3;
        fc1_weights[119][99] = 16'sd-2;
        fc1_weights[119][100] = 16'sd32;
        fc1_weights[119][101] = 16'sd5;
        fc1_weights[119][102] = 16'sd19;
        fc1_weights[119][103] = 16'sd37;
        fc1_weights[119][104] = 16'sd-21;
        fc1_weights[119][105] = 16'sd11;
        fc1_weights[119][106] = 16'sd-17;
        fc1_weights[119][107] = 16'sd-17;
        fc1_weights[119][108] = 16'sd5;
        fc1_weights[119][109] = 16'sd35;
        fc1_weights[119][110] = 16'sd42;
        fc1_weights[119][111] = 16'sd51;
        fc1_weights[119][112] = 16'sd-27;
        fc1_weights[119][113] = 16'sd12;
        fc1_weights[119][114] = 16'sd50;
        fc1_weights[119][115] = 16'sd37;
        fc1_weights[119][116] = 16'sd-1;
        fc1_weights[119][117] = 16'sd23;
        fc1_weights[119][118] = 16'sd56;
        fc1_weights[119][119] = 16'sd8;
        fc1_weights[119][120] = 16'sd5;
        fc1_weights[119][121] = 16'sd-53;
        fc1_weights[119][122] = 16'sd-43;
        fc1_weights[119][123] = 16'sd-26;
        fc1_weights[119][124] = 16'sd14;
        fc1_weights[119][125] = 16'sd6;
        fc1_weights[119][126] = 16'sd41;
        fc1_weights[119][127] = 16'sd-24;
        fc1_weights[119][128] = 16'sd25;
        fc1_weights[119][129] = 16'sd33;
        fc1_weights[119][130] = 16'sd8;
        fc1_weights[119][131] = 16'sd-16;
        fc1_weights[119][132] = 16'sd-14;
        fc1_weights[119][133] = 16'sd-43;
        fc1_weights[119][134] = 16'sd-10;
        fc1_weights[119][135] = 16'sd-5;
        fc1_weights[119][136] = 16'sd16;
        fc1_weights[119][137] = 16'sd41;
        fc1_weights[119][138] = 16'sd-48;
        fc1_weights[119][139] = 16'sd-37;
        fc1_weights[119][140] = 16'sd19;
        fc1_weights[119][141] = 16'sd7;
        fc1_weights[119][142] = 16'sd7;
        fc1_weights[119][143] = 16'sd31;
        fc1_weights[119][144] = 16'sd63;
        fc1_weights[119][145] = 16'sd76;
        fc1_weights[119][146] = 16'sd68;
        fc1_weights[119][147] = 16'sd11;
        fc1_weights[119][148] = 16'sd29;
        fc1_weights[119][149] = 16'sd19;
        fc1_weights[119][150] = 16'sd34;
        fc1_weights[119][151] = 16'sd-33;
        fc1_weights[119][152] = 16'sd10;
        fc1_weights[119][153] = 16'sd-48;
        fc1_weights[119][154] = 16'sd-11;
        fc1_weights[119][155] = 16'sd8;
        fc1_weights[119][156] = 16'sd11;
        fc1_weights[119][157] = 16'sd-3;
        fc1_weights[119][158] = 16'sd39;
        fc1_weights[119][159] = 16'sd24;
        fc1_weights[119][160] = 16'sd30;
        fc1_weights[119][161] = 16'sd32;
        fc1_weights[119][162] = 16'sd2;
        fc1_weights[119][163] = 16'sd-5;
        fc1_weights[119][164] = 16'sd43;
        fc1_weights[119][165] = 16'sd37;
        fc1_weights[119][166] = 16'sd19;
        fc1_weights[119][167] = 16'sd13;
        fc1_weights[119][168] = 16'sd10;
        fc1_weights[119][169] = 16'sd37;
        fc1_weights[119][170] = 16'sd23;
        fc1_weights[119][171] = 16'sd78;
        fc1_weights[119][172] = 16'sd1;
        fc1_weights[119][173] = 16'sd2;
        fc1_weights[119][174] = 16'sd-14;
        fc1_weights[119][175] = 16'sd11;
        fc1_weights[119][176] = 16'sd-26;
        fc1_weights[119][177] = 16'sd-27;
        fc1_weights[119][178] = 16'sd10;
        fc1_weights[119][179] = 16'sd-38;
        fc1_weights[119][180] = 16'sd-39;
        fc1_weights[119][181] = 16'sd-14;
        fc1_weights[119][182] = 16'sd-43;
        fc1_weights[119][183] = 16'sd3;
        fc1_weights[119][184] = 16'sd-11;
        fc1_weights[119][185] = 16'sd2;
        fc1_weights[119][186] = 16'sd23;
        fc1_weights[119][187] = 16'sd6;
        fc1_weights[119][188] = 16'sd12;
        fc1_weights[119][189] = 16'sd9;
        fc1_weights[119][190] = 16'sd-4;
        fc1_weights[119][191] = 16'sd-18;
        fc1_weights[119][192] = 16'sd10;
        fc1_weights[119][193] = 16'sd46;
        fc1_weights[119][194] = 16'sd8;
        fc1_weights[119][195] = 16'sd-10;
        fc1_weights[119][196] = 16'sd7;
        fc1_weights[119][197] = 16'sd0;
        fc1_weights[119][198] = 16'sd38;
        fc1_weights[119][199] = 16'sd17;
        fc1_weights[119][200] = 16'sd-2;
        fc1_weights[119][201] = 16'sd27;
        fc1_weights[119][202] = 16'sd-6;
        fc1_weights[119][203] = 16'sd-86;
        fc1_weights[119][204] = 16'sd-16;
        fc1_weights[119][205] = 16'sd-20;
        fc1_weights[119][206] = 16'sd-6;
        fc1_weights[119][207] = 16'sd-16;
        fc1_weights[120][0] = 16'sd26;
        fc1_weights[120][1] = 16'sd60;
        fc1_weights[120][2] = 16'sd57;
        fc1_weights[120][3] = 16'sd50;
        fc1_weights[120][4] = 16'sd16;
        fc1_weights[120][5] = 16'sd43;
        fc1_weights[120][6] = 16'sd55;
        fc1_weights[120][7] = 16'sd63;
        fc1_weights[120][8] = 16'sd-5;
        fc1_weights[120][9] = 16'sd4;
        fc1_weights[120][10] = 16'sd8;
        fc1_weights[120][11] = 16'sd12;
        fc1_weights[120][12] = 16'sd-19;
        fc1_weights[120][13] = 16'sd-23;
        fc1_weights[120][14] = 16'sd9;
        fc1_weights[120][15] = 16'sd-32;
        fc1_weights[120][16] = 16'sd-4;
        fc1_weights[120][17] = 16'sd-30;
        fc1_weights[120][18] = 16'sd-56;
        fc1_weights[120][19] = 16'sd12;
        fc1_weights[120][20] = 16'sd-34;
        fc1_weights[120][21] = 16'sd29;
        fc1_weights[120][22] = 16'sd12;
        fc1_weights[120][23] = 16'sd29;
        fc1_weights[120][24] = 16'sd-25;
        fc1_weights[120][25] = 16'sd5;
        fc1_weights[120][26] = 16'sd-44;
        fc1_weights[120][27] = 16'sd14;
        fc1_weights[120][28] = 16'sd29;
        fc1_weights[120][29] = 16'sd20;
        fc1_weights[120][30] = 16'sd-14;
        fc1_weights[120][31] = 16'sd-8;
        fc1_weights[120][32] = 16'sd52;
        fc1_weights[120][33] = 16'sd60;
        fc1_weights[120][34] = 16'sd20;
        fc1_weights[120][35] = 16'sd69;
        fc1_weights[120][36] = 16'sd35;
        fc1_weights[120][37] = 16'sd78;
        fc1_weights[120][38] = 16'sd62;
        fc1_weights[120][39] = 16'sd6;
        fc1_weights[120][40] = 16'sd1;
        fc1_weights[120][41] = 16'sd6;
        fc1_weights[120][42] = 16'sd-46;
        fc1_weights[120][43] = 16'sd-12;
        fc1_weights[120][44] = 16'sd18;
        fc1_weights[120][45] = 16'sd27;
        fc1_weights[120][46] = 16'sd10;
        fc1_weights[120][47] = 16'sd-18;
        fc1_weights[120][48] = 16'sd-11;
        fc1_weights[120][49] = 16'sd-25;
        fc1_weights[120][50] = 16'sd50;
        fc1_weights[120][51] = 16'sd29;
        fc1_weights[120][52] = 16'sd-20;
        fc1_weights[120][53] = 16'sd35;
        fc1_weights[120][54] = 16'sd-11;
        fc1_weights[120][55] = 16'sd11;
        fc1_weights[120][56] = 16'sd-14;
        fc1_weights[120][57] = 16'sd-27;
        fc1_weights[120][58] = 16'sd9;
        fc1_weights[120][59] = 16'sd30;
        fc1_weights[120][60] = 16'sd20;
        fc1_weights[120][61] = 16'sd25;
        fc1_weights[120][62] = 16'sd69;
        fc1_weights[120][63] = 16'sd4;
        fc1_weights[120][64] = 16'sd60;
        fc1_weights[120][65] = 16'sd34;
        fc1_weights[120][66] = 16'sd-46;
        fc1_weights[120][67] = 16'sd-32;
        fc1_weights[120][68] = 16'sd19;
        fc1_weights[120][69] = 16'sd38;
        fc1_weights[120][70] = 16'sd41;
        fc1_weights[120][71] = 16'sd-65;
        fc1_weights[120][72] = 16'sd-23;
        fc1_weights[120][73] = 16'sd2;
        fc1_weights[120][74] = 16'sd-21;
        fc1_weights[120][75] = 16'sd-6;
        fc1_weights[120][76] = 16'sd-24;
        fc1_weights[120][77] = 16'sd-5;
        fc1_weights[120][78] = 16'sd-78;
        fc1_weights[120][79] = 16'sd-102;
        fc1_weights[120][80] = 16'sd-20;
        fc1_weights[120][81] = 16'sd-56;
        fc1_weights[120][82] = 16'sd-28;
        fc1_weights[120][83] = 16'sd-19;
        fc1_weights[120][84] = 16'sd2;
        fc1_weights[120][85] = 16'sd14;
        fc1_weights[120][86] = 16'sd20;
        fc1_weights[120][87] = 16'sd-77;
        fc1_weights[120][88] = 16'sd-20;
        fc1_weights[120][89] = 16'sd1;
        fc1_weights[120][90] = 16'sd47;
        fc1_weights[120][91] = 16'sd35;
        fc1_weights[120][92] = 16'sd74;
        fc1_weights[120][93] = 16'sd26;
        fc1_weights[120][94] = 16'sd56;
        fc1_weights[120][95] = 16'sd1;
        fc1_weights[120][96] = 16'sd70;
        fc1_weights[120][97] = 16'sd-26;
        fc1_weights[120][98] = 16'sd-47;
        fc1_weights[120][99] = 16'sd0;
        fc1_weights[120][100] = 16'sd-13;
        fc1_weights[120][101] = 16'sd25;
        fc1_weights[120][102] = 16'sd-6;
        fc1_weights[120][103] = 16'sd-17;
        fc1_weights[120][104] = 16'sd-97;
        fc1_weights[120][105] = 16'sd-10;
        fc1_weights[120][106] = 16'sd-20;
        fc1_weights[120][107] = 16'sd-45;
        fc1_weights[120][108] = 16'sd-85;
        fc1_weights[120][109] = 16'sd-47;
        fc1_weights[120][110] = 16'sd6;
        fc1_weights[120][111] = 16'sd18;
        fc1_weights[120][112] = 16'sd-16;
        fc1_weights[120][113] = 16'sd-66;
        fc1_weights[120][114] = 16'sd-25;
        fc1_weights[120][115] = 16'sd-6;
        fc1_weights[120][116] = 16'sd-39;
        fc1_weights[120][117] = 16'sd5;
        fc1_weights[120][118] = 16'sd8;
        fc1_weights[120][119] = 16'sd-14;
        fc1_weights[120][120] = 16'sd-9;
        fc1_weights[120][121] = 16'sd-1;
        fc1_weights[120][122] = 16'sd28;
        fc1_weights[120][123] = 16'sd-56;
        fc1_weights[120][124] = 16'sd-56;
        fc1_weights[120][125] = 16'sd-11;
        fc1_weights[120][126] = 16'sd-2;
        fc1_weights[120][127] = 16'sd13;
        fc1_weights[120][128] = 16'sd-3;
        fc1_weights[120][129] = 16'sd15;
        fc1_weights[120][130] = 16'sd-20;
        fc1_weights[120][131] = 16'sd-1;
        fc1_weights[120][132] = 16'sd-20;
        fc1_weights[120][133] = 16'sd-34;
        fc1_weights[120][134] = 16'sd-15;
        fc1_weights[120][135] = 16'sd28;
        fc1_weights[120][136] = 16'sd-11;
        fc1_weights[120][137] = 16'sd-48;
        fc1_weights[120][138] = 16'sd37;
        fc1_weights[120][139] = 16'sd63;
        fc1_weights[120][140] = 16'sd-25;
        fc1_weights[120][141] = 16'sd9;
        fc1_weights[120][142] = 16'sd-67;
        fc1_weights[120][143] = 16'sd77;
        fc1_weights[120][144] = 16'sd-28;
        fc1_weights[120][145] = 16'sd24;
        fc1_weights[120][146] = 16'sd33;
        fc1_weights[120][147] = 16'sd4;
        fc1_weights[120][148] = 16'sd-26;
        fc1_weights[120][149] = 16'sd3;
        fc1_weights[120][150] = 16'sd-6;
        fc1_weights[120][151] = 16'sd-6;
        fc1_weights[120][152] = 16'sd10;
        fc1_weights[120][153] = 16'sd8;
        fc1_weights[120][154] = 16'sd-37;
        fc1_weights[120][155] = 16'sd13;
        fc1_weights[120][156] = 16'sd-35;
        fc1_weights[120][157] = 16'sd-43;
        fc1_weights[120][158] = 16'sd-28;
        fc1_weights[120][159] = 16'sd-41;
        fc1_weights[120][160] = 16'sd30;
        fc1_weights[120][161] = 16'sd-17;
        fc1_weights[120][162] = 16'sd7;
        fc1_weights[120][163] = 16'sd14;
        fc1_weights[120][164] = 16'sd4;
        fc1_weights[120][165] = 16'sd-60;
        fc1_weights[120][166] = 16'sd-33;
        fc1_weights[120][167] = 16'sd-35;
        fc1_weights[120][168] = 16'sd-37;
        fc1_weights[120][169] = 16'sd-64;
        fc1_weights[120][170] = 16'sd-65;
        fc1_weights[120][171] = 16'sd-23;
        fc1_weights[120][172] = 16'sd68;
        fc1_weights[120][173] = 16'sd29;
        fc1_weights[120][174] = 16'sd33;
        fc1_weights[120][175] = 16'sd-13;
        fc1_weights[120][176] = 16'sd11;
        fc1_weights[120][177] = 16'sd-36;
        fc1_weights[120][178] = 16'sd-7;
        fc1_weights[120][179] = 16'sd35;
        fc1_weights[120][180] = 16'sd-7;
        fc1_weights[120][181] = 16'sd38;
        fc1_weights[120][182] = 16'sd16;
        fc1_weights[120][183] = 16'sd-2;
        fc1_weights[120][184] = 16'sd11;
        fc1_weights[120][185] = 16'sd11;
        fc1_weights[120][186] = 16'sd66;
        fc1_weights[120][187] = 16'sd60;
        fc1_weights[120][188] = 16'sd44;
        fc1_weights[120][189] = 16'sd35;
        fc1_weights[120][190] = 16'sd-6;
        fc1_weights[120][191] = 16'sd-1;
        fc1_weights[120][192] = 16'sd11;
        fc1_weights[120][193] = 16'sd18;
        fc1_weights[120][194] = 16'sd-38;
        fc1_weights[120][195] = 16'sd-16;
        fc1_weights[120][196] = 16'sd-29;
        fc1_weights[120][197] = 16'sd-39;
        fc1_weights[120][198] = 16'sd6;
        fc1_weights[120][199] = 16'sd24;
        fc1_weights[120][200] = 16'sd44;
        fc1_weights[120][201] = 16'sd11;
        fc1_weights[120][202] = 16'sd-27;
        fc1_weights[120][203] = 16'sd-2;
        fc1_weights[120][204] = 16'sd-7;
        fc1_weights[120][205] = 16'sd38;
        fc1_weights[120][206] = 16'sd7;
        fc1_weights[120][207] = 16'sd9;
        fc1_weights[121][0] = 16'sd3;
        fc1_weights[121][1] = 16'sd5;
        fc1_weights[121][2] = 16'sd43;
        fc1_weights[121][3] = 16'sd-6;
        fc1_weights[121][4] = 16'sd-4;
        fc1_weights[121][5] = 16'sd-4;
        fc1_weights[121][6] = 16'sd-25;
        fc1_weights[121][7] = 16'sd-52;
        fc1_weights[121][8] = 16'sd-7;
        fc1_weights[121][9] = 16'sd29;
        fc1_weights[121][10] = 16'sd59;
        fc1_weights[121][11] = 16'sd82;
        fc1_weights[121][12] = 16'sd19;
        fc1_weights[121][13] = 16'sd40;
        fc1_weights[121][14] = 16'sd4;
        fc1_weights[121][15] = 16'sd-26;
        fc1_weights[121][16] = 16'sd-10;
        fc1_weights[121][17] = 16'sd-3;
        fc1_weights[121][18] = 16'sd-14;
        fc1_weights[121][19] = 16'sd11;
        fc1_weights[121][20] = 16'sd-35;
        fc1_weights[121][21] = 16'sd21;
        fc1_weights[121][22] = 16'sd34;
        fc1_weights[121][23] = 16'sd65;
        fc1_weights[121][24] = 16'sd13;
        fc1_weights[121][25] = 16'sd16;
        fc1_weights[121][26] = 16'sd-8;
        fc1_weights[121][27] = 16'sd14;
        fc1_weights[121][28] = 16'sd24;
        fc1_weights[121][29] = 16'sd46;
        fc1_weights[121][30] = 16'sd31;
        fc1_weights[121][31] = 16'sd84;
        fc1_weights[121][32] = 16'sd-14;
        fc1_weights[121][33] = 16'sd-45;
        fc1_weights[121][34] = 16'sd-41;
        fc1_weights[121][35] = 16'sd-32;
        fc1_weights[121][36] = 16'sd40;
        fc1_weights[121][37] = 16'sd114;
        fc1_weights[121][38] = 16'sd48;
        fc1_weights[121][39] = 16'sd23;
        fc1_weights[121][40] = 16'sd-8;
        fc1_weights[121][41] = 16'sd-42;
        fc1_weights[121][42] = 16'sd-5;
        fc1_weights[121][43] = 16'sd-28;
        fc1_weights[121][44] = 16'sd-20;
        fc1_weights[121][45] = 16'sd-22;
        fc1_weights[121][46] = 16'sd-65;
        fc1_weights[121][47] = 16'sd-29;
        fc1_weights[121][48] = 16'sd-2;
        fc1_weights[121][49] = 16'sd11;
        fc1_weights[121][50] = 16'sd2;
        fc1_weights[121][51] = 16'sd8;
        fc1_weights[121][52] = 16'sd23;
        fc1_weights[121][53] = 16'sd49;
        fc1_weights[121][54] = 16'sd27;
        fc1_weights[121][55] = 16'sd37;
        fc1_weights[121][56] = 16'sd13;
        fc1_weights[121][57] = 16'sd8;
        fc1_weights[121][58] = 16'sd-29;
        fc1_weights[121][59] = 16'sd19;
        fc1_weights[121][60] = 16'sd26;
        fc1_weights[121][61] = 16'sd-37;
        fc1_weights[121][62] = 16'sd-36;
        fc1_weights[121][63] = 16'sd30;
        fc1_weights[121][64] = 16'sd11;
        fc1_weights[121][65] = 16'sd-52;
        fc1_weights[121][66] = 16'sd-13;
        fc1_weights[121][67] = 16'sd-55;
        fc1_weights[121][68] = 16'sd-57;
        fc1_weights[121][69] = 16'sd-11;
        fc1_weights[121][70] = 16'sd2;
        fc1_weights[121][71] = 16'sd-46;
        fc1_weights[121][72] = 16'sd-67;
        fc1_weights[121][73] = 16'sd-36;
        fc1_weights[121][74] = 16'sd-10;
        fc1_weights[121][75] = 16'sd-12;
        fc1_weights[121][76] = 16'sd-1;
        fc1_weights[121][77] = 16'sd-35;
        fc1_weights[121][78] = 16'sd-13;
        fc1_weights[121][79] = 16'sd-53;
        fc1_weights[121][80] = 16'sd47;
        fc1_weights[121][81] = 16'sd43;
        fc1_weights[121][82] = 16'sd-8;
        fc1_weights[121][83] = 16'sd68;
        fc1_weights[121][84] = 16'sd-19;
        fc1_weights[121][85] = 16'sd15;
        fc1_weights[121][86] = 16'sd23;
        fc1_weights[121][87] = 16'sd29;
        fc1_weights[121][88] = 16'sd-15;
        fc1_weights[121][89] = 16'sd-4;
        fc1_weights[121][90] = 16'sd5;
        fc1_weights[121][91] = 16'sd-39;
        fc1_weights[121][92] = 16'sd-34;
        fc1_weights[121][93] = 16'sd20;
        fc1_weights[121][94] = 16'sd-26;
        fc1_weights[121][95] = 16'sd16;
        fc1_weights[121][96] = 16'sd-19;
        fc1_weights[121][97] = 16'sd-12;
        fc1_weights[121][98] = 16'sd-66;
        fc1_weights[121][99] = 16'sd-55;
        fc1_weights[121][100] = 16'sd-12;
        fc1_weights[121][101] = 16'sd-25;
        fc1_weights[121][102] = 16'sd-11;
        fc1_weights[121][103] = 16'sd-4;
        fc1_weights[121][104] = 16'sd34;
        fc1_weights[121][105] = 16'sd5;
        fc1_weights[121][106] = 16'sd41;
        fc1_weights[121][107] = 16'sd30;
        fc1_weights[121][108] = 16'sd30;
        fc1_weights[121][109] = 16'sd48;
        fc1_weights[121][110] = 16'sd-33;
        fc1_weights[121][111] = 16'sd105;
        fc1_weights[121][112] = 16'sd69;
        fc1_weights[121][113] = 16'sd3;
        fc1_weights[121][114] = 16'sd-15;
        fc1_weights[121][115] = 16'sd48;
        fc1_weights[121][116] = 16'sd-73;
        fc1_weights[121][117] = 16'sd1;
        fc1_weights[121][118] = 16'sd-2;
        fc1_weights[121][119] = 16'sd-17;
        fc1_weights[121][120] = 16'sd5;
        fc1_weights[121][121] = 16'sd37;
        fc1_weights[121][122] = 16'sd24;
        fc1_weights[121][123] = 16'sd38;
        fc1_weights[121][124] = 16'sd16;
        fc1_weights[121][125] = 16'sd-21;
        fc1_weights[121][126] = 16'sd42;
        fc1_weights[121][127] = 16'sd33;
        fc1_weights[121][128] = 16'sd17;
        fc1_weights[121][129] = 16'sd9;
        fc1_weights[121][130] = 16'sd-16;
        fc1_weights[121][131] = 16'sd-18;
        fc1_weights[121][132] = 16'sd-41;
        fc1_weights[121][133] = 16'sd-10;
        fc1_weights[121][134] = 16'sd-26;
        fc1_weights[121][135] = 16'sd-30;
        fc1_weights[121][136] = 16'sd2;
        fc1_weights[121][137] = 16'sd21;
        fc1_weights[121][138] = 16'sd7;
        fc1_weights[121][139] = 16'sd-8;
        fc1_weights[121][140] = 16'sd-11;
        fc1_weights[121][141] = 16'sd46;
        fc1_weights[121][142] = 16'sd36;
        fc1_weights[121][143] = 16'sd16;
        fc1_weights[121][144] = 16'sd-10;
        fc1_weights[121][145] = 16'sd31;
        fc1_weights[121][146] = 16'sd-10;
        fc1_weights[121][147] = 16'sd-22;
        fc1_weights[121][148] = 16'sd-12;
        fc1_weights[121][149] = 16'sd-4;
        fc1_weights[121][150] = 16'sd55;
        fc1_weights[121][151] = 16'sd-21;
        fc1_weights[121][152] = 16'sd28;
        fc1_weights[121][153] = 16'sd-65;
        fc1_weights[121][154] = 16'sd8;
        fc1_weights[121][155] = 16'sd2;
        fc1_weights[121][156] = 16'sd-14;
        fc1_weights[121][157] = 16'sd-17;
        fc1_weights[121][158] = 16'sd-32;
        fc1_weights[121][159] = 16'sd-74;
        fc1_weights[121][160] = 16'sd-11;
        fc1_weights[121][161] = 16'sd-8;
        fc1_weights[121][162] = 16'sd52;
        fc1_weights[121][163] = 16'sd15;
        fc1_weights[121][164] = 16'sd-20;
        fc1_weights[121][165] = 16'sd-25;
        fc1_weights[121][166] = 16'sd-22;
        fc1_weights[121][167] = 16'sd-46;
        fc1_weights[121][168] = 16'sd-49;
        fc1_weights[121][169] = 16'sd-53;
        fc1_weights[121][170] = 16'sd-38;
        fc1_weights[121][171] = 16'sd-91;
        fc1_weights[121][172] = 16'sd42;
        fc1_weights[121][173] = 16'sd4;
        fc1_weights[121][174] = 16'sd-20;
        fc1_weights[121][175] = 16'sd-73;
        fc1_weights[121][176] = 16'sd-33;
        fc1_weights[121][177] = 16'sd-39;
        fc1_weights[121][178] = 16'sd-44;
        fc1_weights[121][179] = 16'sd13;
        fc1_weights[121][180] = 16'sd-28;
        fc1_weights[121][181] = 16'sd-1;
        fc1_weights[121][182] = 16'sd-6;
        fc1_weights[121][183] = 16'sd-41;
        fc1_weights[121][184] = 16'sd-35;
        fc1_weights[121][185] = 16'sd8;
        fc1_weights[121][186] = 16'sd108;
        fc1_weights[121][187] = 16'sd20;
        fc1_weights[121][188] = 16'sd31;
        fc1_weights[121][189] = 16'sd51;
        fc1_weights[121][190] = 16'sd1;
        fc1_weights[121][191] = 16'sd-6;
        fc1_weights[121][192] = 16'sd46;
        fc1_weights[121][193] = 16'sd25;
        fc1_weights[121][194] = 16'sd12;
        fc1_weights[121][195] = 16'sd25;
        fc1_weights[121][196] = 16'sd17;
        fc1_weights[121][197] = 16'sd8;
        fc1_weights[121][198] = 16'sd-9;
        fc1_weights[121][199] = 16'sd34;
        fc1_weights[121][200] = 16'sd27;
        fc1_weights[121][201] = 16'sd46;
        fc1_weights[121][202] = 16'sd32;
        fc1_weights[121][203] = 16'sd30;
        fc1_weights[121][204] = 16'sd65;
        fc1_weights[121][205] = 16'sd-15;
        fc1_weights[121][206] = 16'sd-23;
        fc1_weights[121][207] = 16'sd-11;
        fc1_weights[122][0] = 16'sd17;
        fc1_weights[122][1] = 16'sd46;
        fc1_weights[122][2] = 16'sd-34;
        fc1_weights[122][3] = 16'sd-46;
        fc1_weights[122][4] = 16'sd-36;
        fc1_weights[122][5] = 16'sd-1;
        fc1_weights[122][6] = 16'sd-14;
        fc1_weights[122][7] = 16'sd29;
        fc1_weights[122][8] = 16'sd-18;
        fc1_weights[122][9] = 16'sd-55;
        fc1_weights[122][10] = 16'sd65;
        fc1_weights[122][11] = 16'sd7;
        fc1_weights[122][12] = 16'sd-52;
        fc1_weights[122][13] = 16'sd-15;
        fc1_weights[122][14] = 16'sd-96;
        fc1_weights[122][15] = 16'sd18;
        fc1_weights[122][16] = 16'sd-13;
        fc1_weights[122][17] = 16'sd3;
        fc1_weights[122][18] = 16'sd32;
        fc1_weights[122][19] = 16'sd-23;
        fc1_weights[122][20] = 16'sd-14;
        fc1_weights[122][21] = 16'sd2;
        fc1_weights[122][22] = 16'sd-51;
        fc1_weights[122][23] = 16'sd-20;
        fc1_weights[122][24] = 16'sd43;
        fc1_weights[122][25] = 16'sd37;
        fc1_weights[122][26] = 16'sd12;
        fc1_weights[122][27] = 16'sd31;
        fc1_weights[122][28] = 16'sd9;
        fc1_weights[122][29] = 16'sd-13;
        fc1_weights[122][30] = 16'sd-12;
        fc1_weights[122][31] = 16'sd56;
        fc1_weights[122][32] = 16'sd49;
        fc1_weights[122][33] = 16'sd-22;
        fc1_weights[122][34] = 16'sd-29;
        fc1_weights[122][35] = 16'sd-72;
        fc1_weights[122][36] = 16'sd48;
        fc1_weights[122][37] = 16'sd138;
        fc1_weights[122][38] = 16'sd13;
        fc1_weights[122][39] = 16'sd-28;
        fc1_weights[122][40] = 16'sd40;
        fc1_weights[122][41] = 16'sd5;
        fc1_weights[122][42] = 16'sd-38;
        fc1_weights[122][43] = 16'sd51;
        fc1_weights[122][44] = 16'sd25;
        fc1_weights[122][45] = 16'sd28;
        fc1_weights[122][46] = 16'sd6;
        fc1_weights[122][47] = 16'sd-77;
        fc1_weights[122][48] = 16'sd57;
        fc1_weights[122][49] = 16'sd49;
        fc1_weights[122][50] = 16'sd-16;
        fc1_weights[122][51] = 16'sd-39;
        fc1_weights[122][52] = 16'sd7;
        fc1_weights[122][53] = 16'sd49;
        fc1_weights[122][54] = 16'sd-4;
        fc1_weights[122][55] = 16'sd29;
        fc1_weights[122][56] = 16'sd-35;
        fc1_weights[122][57] = 16'sd8;
        fc1_weights[122][58] = 16'sd11;
        fc1_weights[122][59] = 16'sd55;
        fc1_weights[122][60] = 16'sd0;
        fc1_weights[122][61] = 16'sd-31;
        fc1_weights[122][62] = 16'sd-64;
        fc1_weights[122][63] = 16'sd73;
        fc1_weights[122][64] = 16'sd48;
        fc1_weights[122][65] = 16'sd-71;
        fc1_weights[122][66] = 16'sd-47;
        fc1_weights[122][67] = 16'sd-32;
        fc1_weights[122][68] = 16'sd-37;
        fc1_weights[122][69] = 16'sd48;
        fc1_weights[122][70] = 16'sd30;
        fc1_weights[122][71] = 16'sd-17;
        fc1_weights[122][72] = 16'sd-24;
        fc1_weights[122][73] = 16'sd-47;
        fc1_weights[122][74] = 16'sd-50;
        fc1_weights[122][75] = 16'sd-59;
        fc1_weights[122][76] = 16'sd-70;
        fc1_weights[122][77] = 16'sd-43;
        fc1_weights[122][78] = 16'sd18;
        fc1_weights[122][79] = 16'sd33;
        fc1_weights[122][80] = 16'sd-8;
        fc1_weights[122][81] = 16'sd-38;
        fc1_weights[122][82] = 16'sd-40;
        fc1_weights[122][83] = 16'sd4;
        fc1_weights[122][84] = 16'sd24;
        fc1_weights[122][85] = 16'sd-41;
        fc1_weights[122][86] = 16'sd-5;
        fc1_weights[122][87] = 16'sd-36;
        fc1_weights[122][88] = 16'sd6;
        fc1_weights[122][89] = 16'sd28;
        fc1_weights[122][90] = 16'sd14;
        fc1_weights[122][91] = 16'sd-114;
        fc1_weights[122][92] = 16'sd-35;
        fc1_weights[122][93] = 16'sd15;
        fc1_weights[122][94] = 16'sd-79;
        fc1_weights[122][95] = 16'sd48;
        fc1_weights[122][96] = 16'sd-78;
        fc1_weights[122][97] = 16'sd-15;
        fc1_weights[122][98] = 16'sd-25;
        fc1_weights[122][99] = 16'sd-79;
        fc1_weights[122][100] = 16'sd-74;
        fc1_weights[122][101] = 16'sd-61;
        fc1_weights[122][102] = 16'sd-82;
        fc1_weights[122][103] = 16'sd-97;
        fc1_weights[122][104] = 16'sd75;
        fc1_weights[122][105] = 16'sd30;
        fc1_weights[122][106] = 16'sd61;
        fc1_weights[122][107] = 16'sd13;
        fc1_weights[122][108] = 16'sd25;
        fc1_weights[122][109] = 16'sd12;
        fc1_weights[122][110] = 16'sd12;
        fc1_weights[122][111] = 16'sd8;
        fc1_weights[122][112] = 16'sd-12;
        fc1_weights[122][113] = 16'sd57;
        fc1_weights[122][114] = 16'sd67;
        fc1_weights[122][115] = 16'sd59;
        fc1_weights[122][116] = 16'sd-42;
        fc1_weights[122][117] = 16'sd-7;
        fc1_weights[122][118] = 16'sd47;
        fc1_weights[122][119] = 16'sd22;
        fc1_weights[122][120] = 16'sd27;
        fc1_weights[122][121] = 16'sd79;
        fc1_weights[122][122] = 16'sd14;
        fc1_weights[122][123] = 16'sd36;
        fc1_weights[122][124] = 16'sd-26;
        fc1_weights[122][125] = 16'sd-24;
        fc1_weights[122][126] = 16'sd-10;
        fc1_weights[122][127] = 16'sd14;
        fc1_weights[122][128] = 16'sd-32;
        fc1_weights[122][129] = 16'sd-47;
        fc1_weights[122][130] = 16'sd29;
        fc1_weights[122][131] = 16'sd-62;
        fc1_weights[122][132] = 16'sd-33;
        fc1_weights[122][133] = 16'sd-75;
        fc1_weights[122][134] = 16'sd-47;
        fc1_weights[122][135] = 16'sd-44;
        fc1_weights[122][136] = 16'sd-41;
        fc1_weights[122][137] = 16'sd-73;
        fc1_weights[122][138] = 16'sd66;
        fc1_weights[122][139] = 16'sd46;
        fc1_weights[122][140] = 16'sd9;
        fc1_weights[122][141] = 16'sd18;
        fc1_weights[122][142] = 16'sd-7;
        fc1_weights[122][143] = 16'sd54;
        fc1_weights[122][144] = 16'sd29;
        fc1_weights[122][145] = 16'sd28;
        fc1_weights[122][146] = 16'sd60;
        fc1_weights[122][147] = 16'sd37;
        fc1_weights[122][148] = 16'sd-16;
        fc1_weights[122][149] = 16'sd-22;
        fc1_weights[122][150] = 16'sd-16;
        fc1_weights[122][151] = 16'sd-25;
        fc1_weights[122][152] = 16'sd-4;
        fc1_weights[122][153] = 16'sd-41;
        fc1_weights[122][154] = 16'sd-38;
        fc1_weights[122][155] = 16'sd3;
        fc1_weights[122][156] = 16'sd3;
        fc1_weights[122][157] = 16'sd-22;
        fc1_weights[122][158] = 16'sd-44;
        fc1_weights[122][159] = 16'sd5;
        fc1_weights[122][160] = 16'sd8;
        fc1_weights[122][161] = 16'sd-36;
        fc1_weights[122][162] = 16'sd96;
        fc1_weights[122][163] = 16'sd32;
        fc1_weights[122][164] = 16'sd19;
        fc1_weights[122][165] = 16'sd-78;
        fc1_weights[122][166] = 16'sd63;
        fc1_weights[122][167] = 16'sd-14;
        fc1_weights[122][168] = 16'sd0;
        fc1_weights[122][169] = 16'sd-28;
        fc1_weights[122][170] = 16'sd20;
        fc1_weights[122][171] = 16'sd-3;
        fc1_weights[122][172] = 16'sd75;
        fc1_weights[122][173] = 16'sd53;
        fc1_weights[122][174] = 16'sd41;
        fc1_weights[122][175] = 16'sd-3;
        fc1_weights[122][176] = 16'sd29;
        fc1_weights[122][177] = 16'sd36;
        fc1_weights[122][178] = 16'sd-7;
        fc1_weights[122][179] = 16'sd8;
        fc1_weights[122][180] = 16'sd-3;
        fc1_weights[122][181] = 16'sd-4;
        fc1_weights[122][182] = 16'sd30;
        fc1_weights[122][183] = 16'sd22;
        fc1_weights[122][184] = 16'sd-46;
        fc1_weights[122][185] = 16'sd105;
        fc1_weights[122][186] = 16'sd106;
        fc1_weights[122][187] = 16'sd52;
        fc1_weights[122][188] = 16'sd31;
        fc1_weights[122][189] = 16'sd12;
        fc1_weights[122][190] = 16'sd19;
        fc1_weights[122][191] = 16'sd31;
        fc1_weights[122][192] = 16'sd-23;
        fc1_weights[122][193] = 16'sd-41;
        fc1_weights[122][194] = 16'sd-84;
        fc1_weights[122][195] = 16'sd-41;
        fc1_weights[122][196] = 16'sd-11;
        fc1_weights[122][197] = 16'sd-1;
        fc1_weights[122][198] = 16'sd-18;
        fc1_weights[122][199] = 16'sd29;
        fc1_weights[122][200] = 16'sd80;
        fc1_weights[122][201] = 16'sd47;
        fc1_weights[122][202] = 16'sd6;
        fc1_weights[122][203] = 16'sd87;
        fc1_weights[122][204] = 16'sd79;
        fc1_weights[122][205] = 16'sd45;
        fc1_weights[122][206] = 16'sd-10;
        fc1_weights[122][207] = 16'sd28;
        fc1_weights[123][0] = 16'sd18;
        fc1_weights[123][1] = 16'sd-12;
        fc1_weights[123][2] = 16'sd-57;
        fc1_weights[123][3] = 16'sd-15;
        fc1_weights[123][4] = 16'sd-16;
        fc1_weights[123][5] = 16'sd5;
        fc1_weights[123][6] = 16'sd6;
        fc1_weights[123][7] = 16'sd12;
        fc1_weights[123][8] = 16'sd-1;
        fc1_weights[123][9] = 16'sd-8;
        fc1_weights[123][10] = 16'sd-24;
        fc1_weights[123][11] = 16'sd-94;
        fc1_weights[123][12] = 16'sd-111;
        fc1_weights[123][13] = 16'sd19;
        fc1_weights[123][14] = 16'sd90;
        fc1_weights[123][15] = 16'sd79;
        fc1_weights[123][16] = 16'sd77;
        fc1_weights[123][17] = 16'sd-43;
        fc1_weights[123][18] = 16'sd-70;
        fc1_weights[123][19] = 16'sd-82;
        fc1_weights[123][20] = 16'sd20;
        fc1_weights[123][21] = 16'sd-1;
        fc1_weights[123][22] = 16'sd32;
        fc1_weights[123][23] = 16'sd-70;
        fc1_weights[123][24] = 16'sd63;
        fc1_weights[123][25] = 16'sd22;
        fc1_weights[123][26] = 16'sd-20;
        fc1_weights[123][27] = 16'sd-23;
        fc1_weights[123][28] = 16'sd39;
        fc1_weights[123][29] = 16'sd32;
        fc1_weights[123][30] = 16'sd-24;
        fc1_weights[123][31] = 16'sd51;
        fc1_weights[123][32] = 16'sd19;
        fc1_weights[123][33] = 16'sd8;
        fc1_weights[123][34] = 16'sd-32;
        fc1_weights[123][35] = 16'sd-4;
        fc1_weights[123][36] = 16'sd-27;
        fc1_weights[123][37] = 16'sd-98;
        fc1_weights[123][38] = 16'sd-41;
        fc1_weights[123][39] = 16'sd-18;
        fc1_weights[123][40] = 16'sd67;
        fc1_weights[123][41] = 16'sd76;
        fc1_weights[123][42] = 16'sd-4;
        fc1_weights[123][43] = 16'sd-77;
        fc1_weights[123][44] = 16'sd-13;
        fc1_weights[123][45] = 16'sd-74;
        fc1_weights[123][46] = 16'sd2;
        fc1_weights[123][47] = 16'sd-52;
        fc1_weights[123][48] = 16'sd-64;
        fc1_weights[123][49] = 16'sd2;
        fc1_weights[123][50] = 16'sd-1;
        fc1_weights[123][51] = 16'sd-58;
        fc1_weights[123][52] = 16'sd-40;
        fc1_weights[123][53] = 16'sd5;
        fc1_weights[123][54] = 16'sd-46;
        fc1_weights[123][55] = 16'sd-28;
        fc1_weights[123][56] = 16'sd-2;
        fc1_weights[123][57] = 16'sd-24;
        fc1_weights[123][58] = 16'sd40;
        fc1_weights[123][59] = 16'sd-31;
        fc1_weights[123][60] = 16'sd4;
        fc1_weights[123][61] = 16'sd14;
        fc1_weights[123][62] = 16'sd-98;
        fc1_weights[123][63] = 16'sd-23;
        fc1_weights[123][64] = 16'sd-56;
        fc1_weights[123][65] = 16'sd-6;
        fc1_weights[123][66] = 16'sd43;
        fc1_weights[123][67] = 16'sd43;
        fc1_weights[123][68] = 16'sd-24;
        fc1_weights[123][69] = 16'sd-53;
        fc1_weights[123][70] = 16'sd-28;
        fc1_weights[123][71] = 16'sd53;
        fc1_weights[123][72] = 16'sd69;
        fc1_weights[123][73] = 16'sd-4;
        fc1_weights[123][74] = 16'sd-12;
        fc1_weights[123][75] = 16'sd-26;
        fc1_weights[123][76] = 16'sd-39;
        fc1_weights[123][77] = 16'sd14;
        fc1_weights[123][78] = 16'sd32;
        fc1_weights[123][79] = 16'sd132;
        fc1_weights[123][80] = 16'sd27;
        fc1_weights[123][81] = 16'sd-2;
        fc1_weights[123][82] = 16'sd-9;
        fc1_weights[123][83] = 16'sd9;
        fc1_weights[123][84] = 16'sd33;
        fc1_weights[123][85] = 16'sd20;
        fc1_weights[123][86] = 16'sd34;
        fc1_weights[123][87] = 16'sd-21;
        fc1_weights[123][88] = 16'sd-43;
        fc1_weights[123][89] = 16'sd-35;
        fc1_weights[123][90] = 16'sd13;
        fc1_weights[123][91] = 16'sd38;
        fc1_weights[123][92] = 16'sd-16;
        fc1_weights[123][93] = 16'sd43;
        fc1_weights[123][94] = 16'sd0;
        fc1_weights[123][95] = 16'sd22;
        fc1_weights[123][96] = 16'sd-8;
        fc1_weights[123][97] = 16'sd64;
        fc1_weights[123][98] = 16'sd49;
        fc1_weights[123][99] = 16'sd45;
        fc1_weights[123][100] = 16'sd2;
        fc1_weights[123][101] = 16'sd-51;
        fc1_weights[123][102] = 16'sd-13;
        fc1_weights[123][103] = 16'sd2;
        fc1_weights[123][104] = 16'sd62;
        fc1_weights[123][105] = 16'sd-13;
        fc1_weights[123][106] = 16'sd34;
        fc1_weights[123][107] = 16'sd26;
        fc1_weights[123][108] = 16'sd52;
        fc1_weights[123][109] = 16'sd14;
        fc1_weights[123][110] = 16'sd9;
        fc1_weights[123][111] = 16'sd-27;
        fc1_weights[123][112] = 16'sd56;
        fc1_weights[123][113] = 16'sd63;
        fc1_weights[123][114] = 16'sd-26;
        fc1_weights[123][115] = 16'sd-26;
        fc1_weights[123][116] = 16'sd-2;
        fc1_weights[123][117] = 16'sd4;
        fc1_weights[123][118] = 16'sd18;
        fc1_weights[123][119] = 16'sd-23;
        fc1_weights[123][120] = 16'sd-1;
        fc1_weights[123][121] = 16'sd-45;
        fc1_weights[123][122] = 16'sd-26;
        fc1_weights[123][123] = 16'sd-48;
        fc1_weights[123][124] = 16'sd-25;
        fc1_weights[123][125] = 16'sd-31;
        fc1_weights[123][126] = 16'sd-94;
        fc1_weights[123][127] = 16'sd-47;
        fc1_weights[123][128] = 16'sd-47;
        fc1_weights[123][129] = 16'sd-115;
        fc1_weights[123][130] = 16'sd-22;
        fc1_weights[123][131] = 16'sd-36;
        fc1_weights[123][132] = 16'sd3;
        fc1_weights[123][133] = 16'sd-40;
        fc1_weights[123][134] = 16'sd-6;
        fc1_weights[123][135] = 16'sd29;
        fc1_weights[123][136] = 16'sd2;
        fc1_weights[123][137] = 16'sd40;
        fc1_weights[123][138] = 16'sd56;
        fc1_weights[123][139] = 16'sd97;
        fc1_weights[123][140] = 16'sd63;
        fc1_weights[123][141] = 16'sd1;
        fc1_weights[123][142] = 16'sd72;
        fc1_weights[123][143] = 16'sd38;
        fc1_weights[123][144] = 16'sd36;
        fc1_weights[123][145] = 16'sd-6;
        fc1_weights[123][146] = 16'sd-95;
        fc1_weights[123][147] = 16'sd66;
        fc1_weights[123][148] = 16'sd-22;
        fc1_weights[123][149] = 16'sd-75;
        fc1_weights[123][150] = 16'sd-68;
        fc1_weights[123][151] = 16'sd1;
        fc1_weights[123][152] = 16'sd-21;
        fc1_weights[123][153] = 16'sd-15;
        fc1_weights[123][154] = 16'sd14;
        fc1_weights[123][155] = 16'sd54;
        fc1_weights[123][156] = 16'sd-33;
        fc1_weights[123][157] = 16'sd-14;
        fc1_weights[123][158] = 16'sd-6;
        fc1_weights[123][159] = 16'sd5;
        fc1_weights[123][160] = 16'sd-47;
        fc1_weights[123][161] = 16'sd-44;
        fc1_weights[123][162] = 16'sd-24;
        fc1_weights[123][163] = 16'sd38;
        fc1_weights[123][164] = 16'sd-33;
        fc1_weights[123][165] = 16'sd-5;
        fc1_weights[123][166] = 16'sd60;
        fc1_weights[123][167] = 16'sd30;
        fc1_weights[123][168] = 16'sd-48;
        fc1_weights[123][169] = 16'sd5;
        fc1_weights[123][170] = 16'sd52;
        fc1_weights[123][171] = 16'sd4;
        fc1_weights[123][172] = 16'sd-1;
        fc1_weights[123][173] = 16'sd23;
        fc1_weights[123][174] = 16'sd-25;
        fc1_weights[123][175] = 16'sd10;
        fc1_weights[123][176] = 16'sd-7;
        fc1_weights[123][177] = 16'sd-17;
        fc1_weights[123][178] = 16'sd2;
        fc1_weights[123][179] = 16'sd5;
        fc1_weights[123][180] = 16'sd13;
        fc1_weights[123][181] = 16'sd-3;
        fc1_weights[123][182] = 16'sd-3;
        fc1_weights[123][183] = 16'sd-6;
        fc1_weights[123][184] = 16'sd-47;
        fc1_weights[123][185] = 16'sd16;
        fc1_weights[123][186] = 16'sd-46;
        fc1_weights[123][187] = 16'sd-19;
        fc1_weights[123][188] = 16'sd-71;
        fc1_weights[123][189] = 16'sd-34;
        fc1_weights[123][190] = 16'sd4;
        fc1_weights[123][191] = 16'sd18;
        fc1_weights[123][192] = 16'sd40;
        fc1_weights[123][193] = 16'sd36;
        fc1_weights[123][194] = 16'sd42;
        fc1_weights[123][195] = 16'sd26;
        fc1_weights[123][196] = 16'sd14;
        fc1_weights[123][197] = 16'sd28;
        fc1_weights[123][198] = 16'sd2;
        fc1_weights[123][199] = 16'sd44;
        fc1_weights[123][200] = 16'sd-31;
        fc1_weights[123][201] = 16'sd-42;
        fc1_weights[123][202] = 16'sd-38;
        fc1_weights[123][203] = 16'sd66;
        fc1_weights[123][204] = 16'sd-40;
        fc1_weights[123][205] = 16'sd16;
        fc1_weights[123][206] = 16'sd-28;
        fc1_weights[123][207] = 16'sd-22;
        fc1_weights[124][0] = 16'sd-23;
        fc1_weights[124][1] = 16'sd41;
        fc1_weights[124][2] = 16'sd38;
        fc1_weights[124][3] = 16'sd26;
        fc1_weights[124][4] = 16'sd-17;
        fc1_weights[124][5] = 16'sd2;
        fc1_weights[124][6] = 16'sd40;
        fc1_weights[124][7] = 16'sd30;
        fc1_weights[124][8] = 16'sd16;
        fc1_weights[124][9] = 16'sd0;
        fc1_weights[124][10] = 16'sd55;
        fc1_weights[124][11] = 16'sd31;
        fc1_weights[124][12] = 16'sd72;
        fc1_weights[124][13] = 16'sd11;
        fc1_weights[124][14] = 16'sd8;
        fc1_weights[124][15] = 16'sd-16;
        fc1_weights[124][16] = 16'sd-16;
        fc1_weights[124][17] = 16'sd-14;
        fc1_weights[124][18] = 16'sd-31;
        fc1_weights[124][19] = 16'sd-22;
        fc1_weights[124][20] = 16'sd-75;
        fc1_weights[124][21] = 16'sd-11;
        fc1_weights[124][22] = 16'sd-22;
        fc1_weights[124][23] = 16'sd-4;
        fc1_weights[124][24] = 16'sd-51;
        fc1_weights[124][25] = 16'sd-20;
        fc1_weights[124][26] = 16'sd-13;
        fc1_weights[124][27] = 16'sd-3;
        fc1_weights[124][28] = 16'sd8;
        fc1_weights[124][29] = 16'sd33;
        fc1_weights[124][30] = 16'sd3;
        fc1_weights[124][31] = 16'sd-22;
        fc1_weights[124][32] = 16'sd8;
        fc1_weights[124][33] = 16'sd13;
        fc1_weights[124][34] = 16'sd9;
        fc1_weights[124][35] = 16'sd-28;
        fc1_weights[124][36] = 16'sd4;
        fc1_weights[124][37] = 16'sd56;
        fc1_weights[124][38] = 16'sd43;
        fc1_weights[124][39] = 16'sd12;
        fc1_weights[124][40] = 16'sd-3;
        fc1_weights[124][41] = 16'sd-1;
        fc1_weights[124][42] = 16'sd-17;
        fc1_weights[124][43] = 16'sd22;
        fc1_weights[124][44] = 16'sd8;
        fc1_weights[124][45] = 16'sd21;
        fc1_weights[124][46] = 16'sd-35;
        fc1_weights[124][47] = 16'sd-33;
        fc1_weights[124][48] = 16'sd14;
        fc1_weights[124][49] = 16'sd2;
        fc1_weights[124][50] = 16'sd20;
        fc1_weights[124][51] = 16'sd-23;
        fc1_weights[124][52] = 16'sd-27;
        fc1_weights[124][53] = 16'sd29;
        fc1_weights[124][54] = 16'sd1;
        fc1_weights[124][55] = 16'sd43;
        fc1_weights[124][56] = 16'sd8;
        fc1_weights[124][57] = 16'sd-21;
        fc1_weights[124][58] = 16'sd-12;
        fc1_weights[124][59] = 16'sd-2;
        fc1_weights[124][60] = 16'sd-5;
        fc1_weights[124][61] = 16'sd5;
        fc1_weights[124][62] = 16'sd20;
        fc1_weights[124][63] = 16'sd-2;
        fc1_weights[124][64] = 16'sd10;
        fc1_weights[124][65] = 16'sd6;
        fc1_weights[124][66] = 16'sd-27;
        fc1_weights[124][67] = 16'sd-13;
        fc1_weights[124][68] = 16'sd18;
        fc1_weights[124][69] = 16'sd31;
        fc1_weights[124][70] = 16'sd6;
        fc1_weights[124][71] = 16'sd-47;
        fc1_weights[124][72] = 16'sd-52;
        fc1_weights[124][73] = 16'sd6;
        fc1_weights[124][74] = 16'sd22;
        fc1_weights[124][75] = 16'sd3;
        fc1_weights[124][76] = 16'sd-3;
        fc1_weights[124][77] = 16'sd-7;
        fc1_weights[124][78] = 16'sd-51;
        fc1_weights[124][79] = 16'sd-60;
        fc1_weights[124][80] = 16'sd-28;
        fc1_weights[124][81] = 16'sd-1;
        fc1_weights[124][82] = 16'sd17;
        fc1_weights[124][83] = 16'sd-17;
        fc1_weights[124][84] = 16'sd10;
        fc1_weights[124][85] = 16'sd33;
        fc1_weights[124][86] = 16'sd44;
        fc1_weights[124][87] = 16'sd-2;
        fc1_weights[124][88] = 16'sd-18;
        fc1_weights[124][89] = 16'sd9;
        fc1_weights[124][90] = 16'sd-44;
        fc1_weights[124][91] = 16'sd-4;
        fc1_weights[124][92] = 16'sd-8;
        fc1_weights[124][93] = 16'sd-1;
        fc1_weights[124][94] = 16'sd43;
        fc1_weights[124][95] = 16'sd-50;
        fc1_weights[124][96] = 16'sd4;
        fc1_weights[124][97] = 16'sd13;
        fc1_weights[124][98] = 16'sd-44;
        fc1_weights[124][99] = 16'sd2;
        fc1_weights[124][100] = 16'sd-27;
        fc1_weights[124][101] = 16'sd11;
        fc1_weights[124][102] = 16'sd-6;
        fc1_weights[124][103] = 16'sd-7;
        fc1_weights[124][104] = 16'sd-66;
        fc1_weights[124][105] = 16'sd7;
        fc1_weights[124][106] = 16'sd-30;
        fc1_weights[124][107] = 16'sd-17;
        fc1_weights[124][108] = 16'sd22;
        fc1_weights[124][109] = 16'sd7;
        fc1_weights[124][110] = 16'sd-37;
        fc1_weights[124][111] = 16'sd21;
        fc1_weights[124][112] = 16'sd-69;
        fc1_weights[124][113] = 16'sd-64;
        fc1_weights[124][114] = 16'sd-3;
        fc1_weights[124][115] = 16'sd45;
        fc1_weights[124][116] = 16'sd-30;
        fc1_weights[124][117] = 16'sd-50;
        fc1_weights[124][118] = 16'sd-2;
        fc1_weights[124][119] = 16'sd-50;
        fc1_weights[124][120] = 16'sd-55;
        fc1_weights[124][121] = 16'sd-22;
        fc1_weights[124][122] = 16'sd-22;
        fc1_weights[124][123] = 16'sd-37;
        fc1_weights[124][124] = 16'sd-49;
        fc1_weights[124][125] = 16'sd-37;
        fc1_weights[124][126] = 16'sd9;
        fc1_weights[124][127] = 16'sd-27;
        fc1_weights[124][128] = 16'sd-13;
        fc1_weights[124][129] = 16'sd28;
        fc1_weights[124][130] = 16'sd-32;
        fc1_weights[124][131] = 16'sd-5;
        fc1_weights[124][132] = 16'sd-39;
        fc1_weights[124][133] = 16'sd-37;
        fc1_weights[124][134] = 16'sd-2;
        fc1_weights[124][135] = 16'sd2;
        fc1_weights[124][136] = 16'sd18;
        fc1_weights[124][137] = 16'sd-22;
        fc1_weights[124][138] = 16'sd32;
        fc1_weights[124][139] = 16'sd-2;
        fc1_weights[124][140] = 16'sd13;
        fc1_weights[124][141] = 16'sd38;
        fc1_weights[124][142] = 16'sd-6;
        fc1_weights[124][143] = 16'sd68;
        fc1_weights[124][144] = 16'sd40;
        fc1_weights[124][145] = 16'sd41;
        fc1_weights[124][146] = 16'sd20;
        fc1_weights[124][147] = 16'sd-1;
        fc1_weights[124][148] = 16'sd-25;
        fc1_weights[124][149] = 16'sd4;
        fc1_weights[124][150] = 16'sd2;
        fc1_weights[124][151] = 16'sd-39;
        fc1_weights[124][152] = 16'sd16;
        fc1_weights[124][153] = 16'sd-15;
        fc1_weights[124][154] = 16'sd-3;
        fc1_weights[124][155] = 16'sd-37;
        fc1_weights[124][156] = 16'sd-82;
        fc1_weights[124][157] = 16'sd-66;
        fc1_weights[124][158] = 16'sd-23;
        fc1_weights[124][159] = 16'sd-32;
        fc1_weights[124][160] = 16'sd32;
        fc1_weights[124][161] = 16'sd-14;
        fc1_weights[124][162] = 16'sd30;
        fc1_weights[124][163] = 16'sd13;
        fc1_weights[124][164] = 16'sd14;
        fc1_weights[124][165] = 16'sd30;
        fc1_weights[124][166] = 16'sd26;
        fc1_weights[124][167] = 16'sd44;
        fc1_weights[124][168] = 16'sd59;
        fc1_weights[124][169] = 16'sd23;
        fc1_weights[124][170] = 16'sd-3;
        fc1_weights[124][171] = 16'sd34;
        fc1_weights[124][172] = 16'sd47;
        fc1_weights[124][173] = 16'sd18;
        fc1_weights[124][174] = 16'sd13;
        fc1_weights[124][175] = 16'sd-15;
        fc1_weights[124][176] = 16'sd-3;
        fc1_weights[124][177] = 16'sd-12;
        fc1_weights[124][178] = 16'sd-4;
        fc1_weights[124][179] = 16'sd-3;
        fc1_weights[124][180] = 16'sd-18;
        fc1_weights[124][181] = 16'sd13;
        fc1_weights[124][182] = 16'sd-29;
        fc1_weights[124][183] = 16'sd-9;
        fc1_weights[124][184] = 16'sd25;
        fc1_weights[124][185] = 16'sd2;
        fc1_weights[124][186] = 16'sd38;
        fc1_weights[124][187] = 16'sd18;
        fc1_weights[124][188] = 16'sd21;
        fc1_weights[124][189] = 16'sd29;
        fc1_weights[124][190] = 16'sd0;
        fc1_weights[124][191] = 16'sd44;
        fc1_weights[124][192] = 16'sd44;
        fc1_weights[124][193] = 16'sd64;
        fc1_weights[124][194] = 16'sd17;
        fc1_weights[124][195] = 16'sd14;
        fc1_weights[124][196] = 16'sd-4;
        fc1_weights[124][197] = 16'sd-2;
        fc1_weights[124][198] = 16'sd53;
        fc1_weights[124][199] = 16'sd-9;
        fc1_weights[124][200] = 16'sd28;
        fc1_weights[124][201] = 16'sd23;
        fc1_weights[124][202] = 16'sd4;
        fc1_weights[124][203] = 16'sd-3;
        fc1_weights[124][204] = 16'sd33;
        fc1_weights[124][205] = 16'sd-6;
        fc1_weights[124][206] = 16'sd1;
        fc1_weights[124][207] = 16'sd13;
        fc1_weights[125][0] = 16'sd46;
        fc1_weights[125][1] = 16'sd-6;
        fc1_weights[125][2] = 16'sd-20;
        fc1_weights[125][3] = 16'sd-37;
        fc1_weights[125][4] = 16'sd10;
        fc1_weights[125][5] = 16'sd20;
        fc1_weights[125][6] = 16'sd-13;
        fc1_weights[125][7] = 16'sd-59;
        fc1_weights[125][8] = 16'sd-32;
        fc1_weights[125][9] = 16'sd54;
        fc1_weights[125][10] = 16'sd-38;
        fc1_weights[125][11] = 16'sd-4;
        fc1_weights[125][12] = 16'sd-57;
        fc1_weights[125][13] = 16'sd-8;
        fc1_weights[125][14] = 16'sd-44;
        fc1_weights[125][15] = 16'sd3;
        fc1_weights[125][16] = 16'sd-27;
        fc1_weights[125][17] = 16'sd-29;
        fc1_weights[125][18] = 16'sd28;
        fc1_weights[125][19] = 16'sd44;
        fc1_weights[125][20] = 16'sd87;
        fc1_weights[125][21] = 16'sd-25;
        fc1_weights[125][22] = 16'sd9;
        fc1_weights[125][23] = 16'sd30;
        fc1_weights[125][24] = 16'sd49;
        fc1_weights[125][25] = 16'sd-7;
        fc1_weights[125][26] = 16'sd13;
        fc1_weights[125][27] = 16'sd49;
        fc1_weights[125][28] = 16'sd10;
        fc1_weights[125][29] = 16'sd2;
        fc1_weights[125][30] = 16'sd23;
        fc1_weights[125][31] = 16'sd0;
        fc1_weights[125][32] = 16'sd9;
        fc1_weights[125][33] = 16'sd-84;
        fc1_weights[125][34] = 16'sd-79;
        fc1_weights[125][35] = 16'sd-6;
        fc1_weights[125][36] = 16'sd52;
        fc1_weights[125][37] = 16'sd-106;
        fc1_weights[125][38] = 16'sd14;
        fc1_weights[125][39] = 16'sd0;
        fc1_weights[125][40] = 16'sd-5;
        fc1_weights[125][41] = 16'sd-1;
        fc1_weights[125][42] = 16'sd-35;
        fc1_weights[125][43] = 16'sd47;
        fc1_weights[125][44] = 16'sd3;
        fc1_weights[125][45] = 16'sd7;
        fc1_weights[125][46] = 16'sd36;
        fc1_weights[125][47] = 16'sd-19;
        fc1_weights[125][48] = 16'sd6;
        fc1_weights[125][49] = 16'sd8;
        fc1_weights[125][50] = 16'sd-35;
        fc1_weights[125][51] = 16'sd-14;
        fc1_weights[125][52] = 16'sd1;
        fc1_weights[125][53] = 16'sd25;
        fc1_weights[125][54] = 16'sd-4;
        fc1_weights[125][55] = 16'sd19;
        fc1_weights[125][56] = 16'sd34;
        fc1_weights[125][57] = 16'sd41;
        fc1_weights[125][58] = 16'sd-26;
        fc1_weights[125][59] = 16'sd12;
        fc1_weights[125][60] = 16'sd-8;
        fc1_weights[125][61] = 16'sd-19;
        fc1_weights[125][62] = 16'sd-46;
        fc1_weights[125][63] = 16'sd8;
        fc1_weights[125][64] = 16'sd38;
        fc1_weights[125][65] = 16'sd-52;
        fc1_weights[125][66] = 16'sd-49;
        fc1_weights[125][67] = 16'sd1;
        fc1_weights[125][68] = 16'sd-9;
        fc1_weights[125][69] = 16'sd-14;
        fc1_weights[125][70] = 16'sd-26;
        fc1_weights[125][71] = 16'sd19;
        fc1_weights[125][72] = 16'sd1;
        fc1_weights[125][73] = 16'sd-28;
        fc1_weights[125][74] = 16'sd-18;
        fc1_weights[125][75] = 16'sd-14;
        fc1_weights[125][76] = 16'sd32;
        fc1_weights[125][77] = 16'sd-25;
        fc1_weights[125][78] = 16'sd57;
        fc1_weights[125][79] = 16'sd71;
        fc1_weights[125][80] = 16'sd-1;
        fc1_weights[125][81] = 16'sd-30;
        fc1_weights[125][82] = 16'sd-7;
        fc1_weights[125][83] = 16'sd-20;
        fc1_weights[125][84] = 16'sd-13;
        fc1_weights[125][85] = 16'sd-6;
        fc1_weights[125][86] = 16'sd-5;
        fc1_weights[125][87] = 16'sd29;
        fc1_weights[125][88] = 16'sd28;
        fc1_weights[125][89] = 16'sd3;
        fc1_weights[125][90] = 16'sd71;
        fc1_weights[125][91] = 16'sd22;
        fc1_weights[125][92] = 16'sd-16;
        fc1_weights[125][93] = 16'sd-80;
        fc1_weights[125][94] = 16'sd-42;
        fc1_weights[125][95] = 16'sd-6;
        fc1_weights[125][96] = 16'sd-69;
        fc1_weights[125][97] = 16'sd-35;
        fc1_weights[125][98] = 16'sd-6;
        fc1_weights[125][99] = 16'sd-41;
        fc1_weights[125][100] = 16'sd-16;
        fc1_weights[125][101] = 16'sd-42;
        fc1_weights[125][102] = 16'sd-13;
        fc1_weights[125][103] = 16'sd-31;
        fc1_weights[125][104] = 16'sd42;
        fc1_weights[125][105] = 16'sd-5;
        fc1_weights[125][106] = 16'sd7;
        fc1_weights[125][107] = 16'sd44;
        fc1_weights[125][108] = 16'sd47;
        fc1_weights[125][109] = 16'sd20;
        fc1_weights[125][110] = 16'sd42;
        fc1_weights[125][111] = 16'sd-9;
        fc1_weights[125][112] = 16'sd33;
        fc1_weights[125][113] = 16'sd24;
        fc1_weights[125][114] = 16'sd0;
        fc1_weights[125][115] = 16'sd-25;
        fc1_weights[125][116] = 16'sd61;
        fc1_weights[125][117] = 16'sd60;
        fc1_weights[125][118] = 16'sd5;
        fc1_weights[125][119] = 16'sd14;
        fc1_weights[125][120] = 16'sd12;
        fc1_weights[125][121] = 16'sd-3;
        fc1_weights[125][122] = 16'sd-28;
        fc1_weights[125][123] = 16'sd34;
        fc1_weights[125][124] = 16'sd-5;
        fc1_weights[125][125] = 16'sd-2;
        fc1_weights[125][126] = 16'sd-45;
        fc1_weights[125][127] = 16'sd-35;
        fc1_weights[125][128] = 16'sd-50;
        fc1_weights[125][129] = 16'sd-74;
        fc1_weights[125][130] = 16'sd-2;
        fc1_weights[125][131] = 16'sd4;
        fc1_weights[125][132] = 16'sd16;
        fc1_weights[125][133] = 16'sd37;
        fc1_weights[125][134] = 16'sd34;
        fc1_weights[125][135] = 16'sd21;
        fc1_weights[125][136] = 16'sd51;
        fc1_weights[125][137] = 16'sd73;
        fc1_weights[125][138] = 16'sd-6;
        fc1_weights[125][139] = 16'sd10;
        fc1_weights[125][140] = 16'sd-46;
        fc1_weights[125][141] = 16'sd-72;
        fc1_weights[125][142] = 16'sd-20;
        fc1_weights[125][143] = 16'sd-68;
        fc1_weights[125][144] = 16'sd-108;
        fc1_weights[125][145] = 16'sd-111;
        fc1_weights[125][146] = 16'sd-1;
        fc1_weights[125][147] = 16'sd2;
        fc1_weights[125][148] = 16'sd-30;
        fc1_weights[125][149] = 16'sd-47;
        fc1_weights[125][150] = 16'sd-78;
        fc1_weights[125][151] = 16'sd39;
        fc1_weights[125][152] = 16'sd-51;
        fc1_weights[125][153] = 16'sd11;
        fc1_weights[125][154] = 16'sd-63;
        fc1_weights[125][155] = 16'sd65;
        fc1_weights[125][156] = 16'sd27;
        fc1_weights[125][157] = 16'sd24;
        fc1_weights[125][158] = 16'sd-1;
        fc1_weights[125][159] = 16'sd13;
        fc1_weights[125][160] = 16'sd-85;
        fc1_weights[125][161] = 16'sd49;
        fc1_weights[125][162] = 16'sd26;
        fc1_weights[125][163] = 16'sd12;
        fc1_weights[125][164] = 16'sd32;
        fc1_weights[125][165] = 16'sd-44;
        fc1_weights[125][166] = 16'sd-25;
        fc1_weights[125][167] = 16'sd-23;
        fc1_weights[125][168] = 16'sd-77;
        fc1_weights[125][169] = 16'sd9;
        fc1_weights[125][170] = 16'sd-7;
        fc1_weights[125][171] = 16'sd6;
        fc1_weights[125][172] = 16'sd-17;
        fc1_weights[125][173] = 16'sd37;
        fc1_weights[125][174] = 16'sd62;
        fc1_weights[125][175] = 16'sd78;
        fc1_weights[125][176] = 16'sd19;
        fc1_weights[125][177] = 16'sd5;
        fc1_weights[125][178] = 16'sd-1;
        fc1_weights[125][179] = 16'sd20;
        fc1_weights[125][180] = 16'sd-11;
        fc1_weights[125][181] = 16'sd-7;
        fc1_weights[125][182] = 16'sd-46;
        fc1_weights[125][183] = 16'sd-9;
        fc1_weights[125][184] = 16'sd-14;
        fc1_weights[125][185] = 16'sd12;
        fc1_weights[125][186] = 16'sd-15;
        fc1_weights[125][187] = 16'sd0;
        fc1_weights[125][188] = 16'sd-17;
        fc1_weights[125][189] = 16'sd49;
        fc1_weights[125][190] = 16'sd64;
        fc1_weights[125][191] = 16'sd-6;
        fc1_weights[125][192] = 16'sd-47;
        fc1_weights[125][193] = 16'sd-70;
        fc1_weights[125][194] = 16'sd-21;
        fc1_weights[125][195] = 16'sd-25;
        fc1_weights[125][196] = 16'sd38;
        fc1_weights[125][197] = 16'sd46;
        fc1_weights[125][198] = 16'sd10;
        fc1_weights[125][199] = 16'sd2;
        fc1_weights[125][200] = 16'sd15;
        fc1_weights[125][201] = 16'sd13;
        fc1_weights[125][202] = 16'sd-9;
        fc1_weights[125][203] = 16'sd69;
        fc1_weights[125][204] = 16'sd14;
        fc1_weights[125][205] = 16'sd15;
        fc1_weights[125][206] = 16'sd-46;
        fc1_weights[125][207] = 16'sd-58;
        fc1_weights[126][0] = 16'sd-36;
        fc1_weights[126][1] = 16'sd0;
        fc1_weights[126][2] = 16'sd7;
        fc1_weights[126][3] = 16'sd2;
        fc1_weights[126][4] = 16'sd29;
        fc1_weights[126][5] = 16'sd27;
        fc1_weights[126][6] = 16'sd10;
        fc1_weights[126][7] = 16'sd-1;
        fc1_weights[126][8] = 16'sd6;
        fc1_weights[126][9] = 16'sd43;
        fc1_weights[126][10] = 16'sd-4;
        fc1_weights[126][11] = 16'sd-7;
        fc1_weights[126][12] = 16'sd-2;
        fc1_weights[126][13] = 16'sd5;
        fc1_weights[126][14] = 16'sd-29;
        fc1_weights[126][15] = 16'sd-12;
        fc1_weights[126][16] = 16'sd-58;
        fc1_weights[126][17] = 16'sd-63;
        fc1_weights[126][18] = 16'sd-21;
        fc1_weights[126][19] = 16'sd15;
        fc1_weights[126][20] = 16'sd37;
        fc1_weights[126][21] = 16'sd-15;
        fc1_weights[126][22] = 16'sd11;
        fc1_weights[126][23] = 16'sd53;
        fc1_weights[126][24] = 16'sd40;
        fc1_weights[126][25] = 16'sd-33;
        fc1_weights[126][26] = 16'sd8;
        fc1_weights[126][27] = 16'sd9;
        fc1_weights[126][28] = 16'sd3;
        fc1_weights[126][29] = 16'sd-3;
        fc1_weights[126][30] = 16'sd19;
        fc1_weights[126][31] = 16'sd50;
        fc1_weights[126][32] = 16'sd-31;
        fc1_weights[126][33] = 16'sd-40;
        fc1_weights[126][34] = 16'sd-9;
        fc1_weights[126][35] = 16'sd-16;
        fc1_weights[126][36] = 16'sd33;
        fc1_weights[126][37] = 16'sd-24;
        fc1_weights[126][38] = 16'sd7;
        fc1_weights[126][39] = 16'sd0;
        fc1_weights[126][40] = 16'sd-7;
        fc1_weights[126][41] = 16'sd-4;
        fc1_weights[126][42] = 16'sd-43;
        fc1_weights[126][43] = 16'sd-33;
        fc1_weights[126][44] = 16'sd-30;
        fc1_weights[126][45] = 16'sd1;
        fc1_weights[126][46] = 16'sd-16;
        fc1_weights[126][47] = 16'sd-23;
        fc1_weights[126][48] = 16'sd-4;
        fc1_weights[126][49] = 16'sd3;
        fc1_weights[126][50] = 16'sd-2;
        fc1_weights[126][51] = 16'sd-5;
        fc1_weights[126][52] = 16'sd10;
        fc1_weights[126][53] = 16'sd-3;
        fc1_weights[126][54] = 16'sd33;
        fc1_weights[126][55] = 16'sd9;
        fc1_weights[126][56] = 16'sd0;
        fc1_weights[126][57] = 16'sd6;
        fc1_weights[126][58] = 16'sd-27;
        fc1_weights[126][59] = 16'sd-17;
        fc1_weights[126][60] = 16'sd60;
        fc1_weights[126][61] = 16'sd51;
        fc1_weights[126][62] = 16'sd-23;
        fc1_weights[126][63] = 16'sd10;
        fc1_weights[126][64] = 16'sd56;
        fc1_weights[126][65] = 16'sd-47;
        fc1_weights[126][66] = 16'sd-1;
        fc1_weights[126][67] = 16'sd-26;
        fc1_weights[126][68] = 16'sd-38;
        fc1_weights[126][69] = 16'sd-46;
        fc1_weights[126][70] = 16'sd-26;
        fc1_weights[126][71] = 16'sd35;
        fc1_weights[126][72] = 16'sd3;
        fc1_weights[126][73] = 16'sd-5;
        fc1_weights[126][74] = 16'sd-17;
        fc1_weights[126][75] = 16'sd3;
        fc1_weights[126][76] = 16'sd12;
        fc1_weights[126][77] = 16'sd-17;
        fc1_weights[126][78] = 16'sd-8;
        fc1_weights[126][79] = 16'sd51;
        fc1_weights[126][80] = 16'sd8;
        fc1_weights[126][81] = 16'sd51;
        fc1_weights[126][82] = 16'sd9;
        fc1_weights[126][83] = 16'sd38;
        fc1_weights[126][84] = 16'sd-24;
        fc1_weights[126][85] = 16'sd-16;
        fc1_weights[126][86] = 16'sd64;
        fc1_weights[126][87] = 16'sd99;
        fc1_weights[126][88] = 16'sd53;
        fc1_weights[126][89] = 16'sd49;
        fc1_weights[126][90] = 16'sd124;
        fc1_weights[126][91] = 16'sd65;
        fc1_weights[126][92] = 16'sd-27;
        fc1_weights[126][93] = 16'sd-58;
        fc1_weights[126][94] = 16'sd-74;
        fc1_weights[126][95] = 16'sd-38;
        fc1_weights[126][96] = 16'sd-13;
        fc1_weights[126][97] = 16'sd-12;
        fc1_weights[126][98] = 16'sd10;
        fc1_weights[126][99] = 16'sd-35;
        fc1_weights[126][100] = 16'sd4;
        fc1_weights[126][101] = 16'sd-34;
        fc1_weights[126][102] = 16'sd-12;
        fc1_weights[126][103] = 16'sd-16;
        fc1_weights[126][104] = 16'sd-4;
        fc1_weights[126][105] = 16'sd-29;
        fc1_weights[126][106] = 16'sd4;
        fc1_weights[126][107] = 16'sd36;
        fc1_weights[126][108] = 16'sd30;
        fc1_weights[126][109] = 16'sd39;
        fc1_weights[126][110] = 16'sd8;
        fc1_weights[126][111] = 16'sd12;
        fc1_weights[126][112] = 16'sd62;
        fc1_weights[126][113] = 16'sd47;
        fc1_weights[126][114] = 16'sd39;
        fc1_weights[126][115] = 16'sd36;
        fc1_weights[126][116] = 16'sd64;
        fc1_weights[126][117] = 16'sd78;
        fc1_weights[126][118] = 16'sd-2;
        fc1_weights[126][119] = 16'sd-2;
        fc1_weights[126][120] = 16'sd2;
        fc1_weights[126][121] = 16'sd-11;
        fc1_weights[126][122] = 16'sd-4;
        fc1_weights[126][123] = 16'sd12;
        fc1_weights[126][124] = 16'sd-8;
        fc1_weights[126][125] = 16'sd-20;
        fc1_weights[126][126] = 16'sd-19;
        fc1_weights[126][127] = 16'sd-4;
        fc1_weights[126][128] = 16'sd-20;
        fc1_weights[126][129] = 16'sd-43;
        fc1_weights[126][130] = 16'sd21;
        fc1_weights[126][131] = 16'sd23;
        fc1_weights[126][132] = 16'sd48;
        fc1_weights[126][133] = 16'sd45;
        fc1_weights[126][134] = 16'sd-3;
        fc1_weights[126][135] = 16'sd42;
        fc1_weights[126][136] = 16'sd12;
        fc1_weights[126][137] = 16'sd54;
        fc1_weights[126][138] = 16'sd3;
        fc1_weights[126][139] = 16'sd-5;
        fc1_weights[126][140] = 16'sd-38;
        fc1_weights[126][141] = 16'sd-35;
        fc1_weights[126][142] = 16'sd48;
        fc1_weights[126][143] = 16'sd7;
        fc1_weights[126][144] = 16'sd-14;
        fc1_weights[126][145] = 16'sd-47;
        fc1_weights[126][146] = 16'sd-2;
        fc1_weights[126][147] = 16'sd-27;
        fc1_weights[126][148] = 16'sd-2;
        fc1_weights[126][149] = 16'sd-38;
        fc1_weights[126][150] = 16'sd-34;
        fc1_weights[126][151] = 16'sd-16;
        fc1_weights[126][152] = 16'sd-34;
        fc1_weights[126][153] = 16'sd-47;
        fc1_weights[126][154] = 16'sd-44;
        fc1_weights[126][155] = 16'sd-9;
        fc1_weights[126][156] = 16'sd11;
        fc1_weights[126][157] = 16'sd12;
        fc1_weights[126][158] = 16'sd-12;
        fc1_weights[126][159] = 16'sd-1;
        fc1_weights[126][160] = 16'sd-62;
        fc1_weights[126][161] = 16'sd5;
        fc1_weights[126][162] = 16'sd1;
        fc1_weights[126][163] = 16'sd6;
        fc1_weights[126][164] = 16'sd-1;
        fc1_weights[126][165] = 16'sd-64;
        fc1_weights[126][166] = 16'sd-39;
        fc1_weights[126][167] = 16'sd-25;
        fc1_weights[126][168] = 16'sd-16;
        fc1_weights[126][169] = 16'sd3;
        fc1_weights[126][170] = 16'sd-7;
        fc1_weights[126][171] = 16'sd-1;
        fc1_weights[126][172] = 16'sd-6;
        fc1_weights[126][173] = 16'sd-24;
        fc1_weights[126][174] = 16'sd12;
        fc1_weights[126][175] = 16'sd38;
        fc1_weights[126][176] = 16'sd12;
        fc1_weights[126][177] = 16'sd-40;
        fc1_weights[126][178] = 16'sd-5;
        fc1_weights[126][179] = 16'sd10;
        fc1_weights[126][180] = 16'sd-11;
        fc1_weights[126][181] = 16'sd-27;
        fc1_weights[126][182] = 16'sd-5;
        fc1_weights[126][183] = 16'sd-7;
        fc1_weights[126][184] = 16'sd-15;
        fc1_weights[126][185] = 16'sd-27;
        fc1_weights[126][186] = 16'sd-89;
        fc1_weights[126][187] = 16'sd-53;
        fc1_weights[126][188] = 16'sd-32;
        fc1_weights[126][189] = 16'sd5;
        fc1_weights[126][190] = 16'sd7;
        fc1_weights[126][191] = 16'sd-7;
        fc1_weights[126][192] = 16'sd-16;
        fc1_weights[126][193] = 16'sd-27;
        fc1_weights[126][194] = 16'sd-6;
        fc1_weights[126][195] = 16'sd-17;
        fc1_weights[126][196] = 16'sd-7;
        fc1_weights[126][197] = 16'sd31;
        fc1_weights[126][198] = 16'sd-19;
        fc1_weights[126][199] = 16'sd-6;
        fc1_weights[126][200] = 16'sd8;
        fc1_weights[126][201] = 16'sd20;
        fc1_weights[126][202] = 16'sd-7;
        fc1_weights[126][203] = 16'sd46;
        fc1_weights[126][204] = 16'sd26;
        fc1_weights[126][205] = 16'sd-20;
        fc1_weights[126][206] = 16'sd-50;
        fc1_weights[126][207] = 16'sd-38;
        fc1_weights[127][0] = 16'sd-4;
        fc1_weights[127][1] = 16'sd-2;
        fc1_weights[127][2] = 16'sd40;
        fc1_weights[127][3] = 16'sd14;
        fc1_weights[127][4] = 16'sd14;
        fc1_weights[127][5] = 16'sd22;
        fc1_weights[127][6] = 16'sd35;
        fc1_weights[127][7] = 16'sd1;
        fc1_weights[127][8] = 16'sd6;
        fc1_weights[127][9] = 16'sd58;
        fc1_weights[127][10] = 16'sd41;
        fc1_weights[127][11] = 16'sd0;
        fc1_weights[127][12] = 16'sd-3;
        fc1_weights[127][13] = 16'sd-4;
        fc1_weights[127][14] = 16'sd-16;
        fc1_weights[127][15] = 16'sd30;
        fc1_weights[127][16] = 16'sd-20;
        fc1_weights[127][17] = 16'sd2;
        fc1_weights[127][18] = 16'sd36;
        fc1_weights[127][19] = 16'sd-17;
        fc1_weights[127][20] = 16'sd-14;
        fc1_weights[127][21] = 16'sd-38;
        fc1_weights[127][22] = 16'sd25;
        fc1_weights[127][23] = 16'sd4;
        fc1_weights[127][24] = 16'sd41;
        fc1_weights[127][25] = 16'sd28;
        fc1_weights[127][26] = 16'sd-62;
        fc1_weights[127][27] = 16'sd7;
        fc1_weights[127][28] = 16'sd12;
        fc1_weights[127][29] = 16'sd17;
        fc1_weights[127][30] = 16'sd16;
        fc1_weights[127][31] = 16'sd59;
        fc1_weights[127][32] = 16'sd27;
        fc1_weights[127][33] = 16'sd-41;
        fc1_weights[127][34] = 16'sd13;
        fc1_weights[127][35] = 16'sd5;
        fc1_weights[127][36] = 16'sd26;
        fc1_weights[127][37] = 16'sd50;
        fc1_weights[127][38] = 16'sd-46;
        fc1_weights[127][39] = 16'sd-62;
        fc1_weights[127][40] = 16'sd46;
        fc1_weights[127][41] = 16'sd25;
        fc1_weights[127][42] = 16'sd7;
        fc1_weights[127][43] = 16'sd57;
        fc1_weights[127][44] = 16'sd54;
        fc1_weights[127][45] = 16'sd34;
        fc1_weights[127][46] = 16'sd-43;
        fc1_weights[127][47] = 16'sd2;
        fc1_weights[127][48] = 16'sd-17;
        fc1_weights[127][49] = 16'sd48;
        fc1_weights[127][50] = 16'sd-15;
        fc1_weights[127][51] = 16'sd1;
        fc1_weights[127][52] = 16'sd-36;
        fc1_weights[127][53] = 16'sd-48;
        fc1_weights[127][54] = 16'sd-11;
        fc1_weights[127][55] = 16'sd-59;
        fc1_weights[127][56] = 16'sd-10;
        fc1_weights[127][57] = 16'sd-16;
        fc1_weights[127][58] = 16'sd-64;
        fc1_weights[127][59] = 16'sd-49;
        fc1_weights[127][60] = 16'sd-15;
        fc1_weights[127][61] = 16'sd-74;
        fc1_weights[127][62] = 16'sd23;
        fc1_weights[127][63] = 16'sd39;
        fc1_weights[127][64] = 16'sd-59;
        fc1_weights[127][65] = 16'sd-18;
        fc1_weights[127][66] = 16'sd-3;
        fc1_weights[127][67] = 16'sd-11;
        fc1_weights[127][68] = 16'sd20;
        fc1_weights[127][69] = 16'sd-3;
        fc1_weights[127][70] = 16'sd31;
        fc1_weights[127][71] = 16'sd-45;
        fc1_weights[127][72] = 16'sd-35;
        fc1_weights[127][73] = 16'sd2;
        fc1_weights[127][74] = 16'sd6;
        fc1_weights[127][75] = 16'sd23;
        fc1_weights[127][76] = 16'sd59;
        fc1_weights[127][77] = 16'sd-4;
        fc1_weights[127][78] = 16'sd-14;
        fc1_weights[127][79] = 16'sd-2;
        fc1_weights[127][80] = 16'sd8;
        fc1_weights[127][81] = 16'sd-46;
        fc1_weights[127][82] = 16'sd-10;
        fc1_weights[127][83] = 16'sd-60;
        fc1_weights[127][84] = 16'sd-64;
        fc1_weights[127][85] = 16'sd-69;
        fc1_weights[127][86] = 16'sd-79;
        fc1_weights[127][87] = 16'sd-32;
        fc1_weights[127][88] = 16'sd-61;
        fc1_weights[127][89] = 16'sd41;
        fc1_weights[127][90] = 16'sd-32;
        fc1_weights[127][91] = 16'sd-29;
        fc1_weights[127][92] = 16'sd-49;
        fc1_weights[127][93] = 16'sd25;
        fc1_weights[127][94] = 16'sd-26;
        fc1_weights[127][95] = 16'sd7;
        fc1_weights[127][96] = 16'sd13;
        fc1_weights[127][97] = 16'sd-22;
        fc1_weights[127][98] = 16'sd-27;
        fc1_weights[127][99] = 16'sd-14;
        fc1_weights[127][100] = 16'sd42;
        fc1_weights[127][101] = 16'sd46;
        fc1_weights[127][102] = 16'sd34;
        fc1_weights[127][103] = 16'sd-8;
        fc1_weights[127][104] = 16'sd-25;
        fc1_weights[127][105] = 16'sd13;
        fc1_weights[127][106] = 16'sd-19;
        fc1_weights[127][107] = 16'sd-18;
        fc1_weights[127][108] = 16'sd6;
        fc1_weights[127][109] = 16'sd-19;
        fc1_weights[127][110] = 16'sd-5;
        fc1_weights[127][111] = 16'sd6;
        fc1_weights[127][112] = 16'sd10;
        fc1_weights[127][113] = 16'sd-2;
        fc1_weights[127][114] = 16'sd-4;
        fc1_weights[127][115] = 16'sd-34;
        fc1_weights[127][116] = 16'sd1;
        fc1_weights[127][117] = 16'sd31;
        fc1_weights[127][118] = 16'sd27;
        fc1_weights[127][119] = 16'sd102;
        fc1_weights[127][120] = 16'sd23;
        fc1_weights[127][121] = 16'sd56;
        fc1_weights[127][122] = 16'sd66;
        fc1_weights[127][123] = 16'sd18;
        fc1_weights[127][124] = 16'sd33;
        fc1_weights[127][125] = 16'sd26;
        fc1_weights[127][126] = 16'sd18;
        fc1_weights[127][127] = 16'sd13;
        fc1_weights[127][128] = 16'sd10;
        fc1_weights[127][129] = 16'sd-2;
        fc1_weights[127][130] = 16'sd-3;
        fc1_weights[127][131] = 16'sd13;
        fc1_weights[127][132] = 16'sd42;
        fc1_weights[127][133] = 16'sd-12;
        fc1_weights[127][134] = 16'sd-3;
        fc1_weights[127][135] = 16'sd-6;
        fc1_weights[127][136] = 16'sd-40;
        fc1_weights[127][137] = 16'sd13;
        fc1_weights[127][138] = 16'sd-27;
        fc1_weights[127][139] = 16'sd18;
        fc1_weights[127][140] = 16'sd16;
        fc1_weights[127][141] = 16'sd-1;
        fc1_weights[127][142] = 16'sd94;
        fc1_weights[127][143] = 16'sd16;
        fc1_weights[127][144] = 16'sd-1;
        fc1_weights[127][145] = 16'sd-44;
        fc1_weights[127][146] = 16'sd8;
        fc1_weights[127][147] = 16'sd-28;
        fc1_weights[127][148] = 16'sd23;
        fc1_weights[127][149] = 16'sd25;
        fc1_weights[127][150] = 16'sd46;
        fc1_weights[127][151] = 16'sd-22;
        fc1_weights[127][152] = 16'sd-12;
        fc1_weights[127][153] = 16'sd4;
        fc1_weights[127][154] = 16'sd1;
        fc1_weights[127][155] = 16'sd-7;
        fc1_weights[127][156] = 16'sd35;
        fc1_weights[127][157] = 16'sd43;
        fc1_weights[127][158] = 16'sd5;
        fc1_weights[127][159] = 16'sd-20;
        fc1_weights[127][160] = 16'sd-32;
        fc1_weights[127][161] = 16'sd-46;
        fc1_weights[127][162] = 16'sd7;
        fc1_weights[127][163] = 16'sd-29;
        fc1_weights[127][164] = 16'sd-11;
        fc1_weights[127][165] = 16'sd13;
        fc1_weights[127][166] = 16'sd28;
        fc1_weights[127][167] = 16'sd18;
        fc1_weights[127][168] = 16'sd83;
        fc1_weights[127][169] = 16'sd40;
        fc1_weights[127][170] = 16'sd28;
        fc1_weights[127][171] = 16'sd37;
        fc1_weights[127][172] = 16'sd40;
        fc1_weights[127][173] = 16'sd62;
        fc1_weights[127][174] = 16'sd42;
        fc1_weights[127][175] = 16'sd18;
        fc1_weights[127][176] = 16'sd27;
        fc1_weights[127][177] = 16'sd47;
        fc1_weights[127][178] = 16'sd6;
        fc1_weights[127][179] = 16'sd53;
        fc1_weights[127][180] = 16'sd26;
        fc1_weights[127][181] = 16'sd0;
        fc1_weights[127][182] = 16'sd40;
        fc1_weights[127][183] = 16'sd20;
        fc1_weights[127][184] = 16'sd13;
        fc1_weights[127][185] = 16'sd21;
        fc1_weights[127][186] = 16'sd22;
        fc1_weights[127][187] = 16'sd31;
        fc1_weights[127][188] = 16'sd1;
        fc1_weights[127][189] = 16'sd-15;
        fc1_weights[127][190] = 16'sd11;
        fc1_weights[127][191] = 16'sd7;
        fc1_weights[127][192] = 16'sd-27;
        fc1_weights[127][193] = 16'sd-9;
        fc1_weights[127][194] = 16'sd46;
        fc1_weights[127][195] = 16'sd47;
        fc1_weights[127][196] = 16'sd12;
        fc1_weights[127][197] = 16'sd30;
        fc1_weights[127][198] = 16'sd16;
        fc1_weights[127][199] = 16'sd25;
        fc1_weights[127][200] = 16'sd1;
        fc1_weights[127][201] = 16'sd20;
        fc1_weights[127][202] = 16'sd41;
        fc1_weights[127][203] = 16'sd35;
        fc1_weights[127][204] = 16'sd32;
        fc1_weights[127][205] = 16'sd42;
        fc1_weights[127][206] = 16'sd26;
        fc1_weights[127][207] = 16'sd-16;
        // fc1 biases
        fc1_biases[0] = 16'sd0;
        fc1_biases[1] = 16'sd0;
        fc1_biases[2] = 16'sd0;
        fc1_biases[3] = 16'sd0;
        fc1_biases[4] = 16'sd0;
        fc1_biases[5] = 16'sd0;
        fc1_biases[6] = 16'sd0;
        fc1_biases[7] = 16'sd0;
        fc1_biases[8] = 16'sd0;
        fc1_biases[9] = 16'sd0;
        fc1_biases[10] = 16'sd0;
        fc1_biases[11] = 16'sd0;
        fc1_biases[12] = 16'sd0;
        fc1_biases[13] = 16'sd0;
        fc1_biases[14] = 16'sd0;
        fc1_biases[15] = 16'sd0;
        fc1_biases[16] = 16'sd0;
        fc1_biases[17] = 16'sd0;
        fc1_biases[18] = 16'sd0;
        fc1_biases[19] = 16'sd0;
        fc1_biases[20] = 16'sd0;
        fc1_biases[21] = 16'sd0;
        fc1_biases[22] = 16'sd0;
        fc1_biases[23] = 16'sd0;
        fc1_biases[24] = 16'sd0;
        fc1_biases[25] = 16'sd0;
        fc1_biases[26] = 16'sd0;
        fc1_biases[27] = 16'sd0;
        fc1_biases[28] = 16'sd0;
        fc1_biases[29] = 16'sd0;
        fc1_biases[30] = 16'sd0;
        fc1_biases[31] = 16'sd0;
        fc1_biases[32] = 16'sd0;
        fc1_biases[33] = 16'sd0;
        fc1_biases[34] = 16'sd0;
        fc1_biases[35] = 16'sd0;
        fc1_biases[36] = 16'sd0;
        fc1_biases[37] = 16'sd0;
        fc1_biases[38] = 16'sd0;
        fc1_biases[39] = 16'sd0;
        fc1_biases[40] = 16'sd0;
        fc1_biases[41] = 16'sd0;
        fc1_biases[42] = 16'sd0;
        fc1_biases[43] = 16'sd0;
        fc1_biases[44] = 16'sd0;
        fc1_biases[45] = 16'sd0;
        fc1_biases[46] = 16'sd0;
        fc1_biases[47] = 16'sd0;
        fc1_biases[48] = 16'sd0;
        fc1_biases[49] = 16'sd0;
        fc1_biases[50] = 16'sd0;
        fc1_biases[51] = 16'sd0;
        fc1_biases[52] = 16'sd0;
        fc1_biases[53] = 16'sd0;
        fc1_biases[54] = 16'sd0;
        fc1_biases[55] = 16'sd0;
        fc1_biases[56] = 16'sd0;
        fc1_biases[57] = 16'sd0;
        fc1_biases[58] = 16'sd0;
        fc1_biases[59] = 16'sd0;
        fc1_biases[60] = 16'sd0;
        fc1_biases[61] = 16'sd0;
        fc1_biases[62] = 16'sd0;
        fc1_biases[63] = 16'sd0;
        fc1_biases[64] = 16'sd0;
        fc1_biases[65] = 16'sd0;
        fc1_biases[66] = 16'sd0;
        fc1_biases[67] = 16'sd0;
        fc1_biases[68] = 16'sd0;
        fc1_biases[69] = 16'sd0;
        fc1_biases[70] = 16'sd0;
        fc1_biases[71] = 16'sd0;
        fc1_biases[72] = 16'sd0;
        fc1_biases[73] = 16'sd0;
        fc1_biases[74] = 16'sd0;
        fc1_biases[75] = 16'sd0;
        fc1_biases[76] = 16'sd0;
        fc1_biases[77] = 16'sd0;
        fc1_biases[78] = 16'sd0;
        fc1_biases[79] = 16'sd0;
        fc1_biases[80] = 16'sd0;
        fc1_biases[81] = 16'sd0;
        fc1_biases[82] = 16'sd0;
        fc1_biases[83] = 16'sd0;
        fc1_biases[84] = 16'sd0;
        fc1_biases[85] = 16'sd0;
        fc1_biases[86] = 16'sd0;
        fc1_biases[87] = 16'sd0;
        fc1_biases[88] = 16'sd0;
        fc1_biases[89] = 16'sd0;
        fc1_biases[90] = 16'sd0;
        fc1_biases[91] = 16'sd0;
        fc1_biases[92] = 16'sd0;
        fc1_biases[93] = 16'sd0;
        fc1_biases[94] = 16'sd0;
        fc1_biases[95] = 16'sd0;
        fc1_biases[96] = 16'sd0;
        fc1_biases[97] = 16'sd0;
        fc1_biases[98] = 16'sd0;
        fc1_biases[99] = 16'sd0;
        fc1_biases[100] = 16'sd0;
        fc1_biases[101] = 16'sd0;
        fc1_biases[102] = 16'sd0;
        fc1_biases[103] = 16'sd0;
        fc1_biases[104] = 16'sd0;
        fc1_biases[105] = 16'sd0;
        fc1_biases[106] = 16'sd0;
        fc1_biases[107] = 16'sd0;
        fc1_biases[108] = 16'sd0;
        fc1_biases[109] = 16'sd0;
        fc1_biases[110] = 16'sd0;
        fc1_biases[111] = 16'sd0;
        fc1_biases[112] = 16'sd0;
        fc1_biases[113] = 16'sd0;
        fc1_biases[114] = 16'sd0;
        fc1_biases[115] = 16'sd0;
        fc1_biases[116] = 16'sd0;
        fc1_biases[117] = 16'sd0;
        fc1_biases[118] = 16'sd0;
        fc1_biases[119] = 16'sd0;
        fc1_biases[120] = 16'sd0;
        fc1_biases[121] = 16'sd0;
        fc1_biases[122] = 16'sd0;
        fc1_biases[123] = 16'sd0;
        fc1_biases[124] = 16'sd0;
        fc1_biases[125] = 16'sd0;
        fc1_biases[126] = 16'sd0;
        fc1_biases[127] = 16'sd0;
        
        // fc2 weights
        fc2_weights[0][0] = 16'sd-11;
        fc2_weights[0][1] = 16'sd-28;
        fc2_weights[0][2] = 16'sd3;
        fc2_weights[0][3] = 16'sd60;
        fc2_weights[0][4] = 16'sd-49;
        fc2_weights[0][5] = 16'sd39;
        fc2_weights[0][6] = 16'sd-60;
        fc2_weights[0][7] = 16'sd-45;
        fc2_weights[0][8] = 16'sd-52;
        fc2_weights[0][9] = 16'sd1;
        fc2_weights[0][10] = 16'sd-44;
        fc2_weights[0][11] = 16'sd-58;
        fc2_weights[0][12] = 16'sd38;
        fc2_weights[0][13] = 16'sd49;
        fc2_weights[0][14] = 16'sd17;
        fc2_weights[0][15] = 16'sd60;
        fc2_weights[0][16] = 16'sd-14;
        fc2_weights[0][17] = 16'sd-4;
        fc2_weights[0][18] = 16'sd-33;
        fc2_weights[0][19] = 16'sd28;
        fc2_weights[0][20] = 16'sd40;
        fc2_weights[0][21] = 16'sd-34;
        fc2_weights[0][22] = 16'sd-39;
        fc2_weights[0][23] = 16'sd-42;
        fc2_weights[0][24] = 16'sd9;
        fc2_weights[0][25] = 16'sd27;
        fc2_weights[0][26] = 16'sd11;
        fc2_weights[0][27] = 16'sd35;
        fc2_weights[0][28] = 16'sd-23;
        fc2_weights[0][29] = 16'sd-52;
        fc2_weights[0][30] = 16'sd24;
        fc2_weights[0][31] = 16'sd-52;
        fc2_weights[0][32] = 16'sd12;
        fc2_weights[0][33] = 16'sd4;
        fc2_weights[0][34] = 16'sd21;
        fc2_weights[0][35] = 16'sd47;
        fc2_weights[0][36] = 16'sd-27;
        fc2_weights[0][37] = 16'sd0;
        fc2_weights[0][38] = 16'sd-60;
        fc2_weights[0][39] = 16'sd-19;
        fc2_weights[0][40] = 16'sd37;
        fc2_weights[0][41] = 16'sd0;
        fc2_weights[0][42] = 16'sd13;
        fc2_weights[0][43] = 16'sd-19;
        fc2_weights[0][44] = 16'sd61;
        fc2_weights[0][45] = 16'sd61;
        fc2_weights[0][46] = 16'sd0;
        fc2_weights[0][47] = 16'sd25;
        fc2_weights[0][48] = 16'sd30;
        fc2_weights[0][49] = 16'sd-15;
        fc2_weights[0][50] = 16'sd37;
        fc2_weights[0][51] = 16'sd2;
        fc2_weights[0][52] = 16'sd-7;
        fc2_weights[0][53] = 16'sd-18;
        fc2_weights[0][54] = 16'sd-30;
        fc2_weights[0][55] = 16'sd-14;
        fc2_weights[0][56] = 16'sd9;
        fc2_weights[0][57] = 16'sd12;
        fc2_weights[0][58] = 16'sd54;
        fc2_weights[0][59] = 16'sd19;
        fc2_weights[0][60] = 16'sd-40;
        fc2_weights[0][61] = 16'sd-41;
        fc2_weights[0][62] = 16'sd32;
        fc2_weights[0][63] = 16'sd42;
        fc2_weights[0][64] = 16'sd-88;
        fc2_weights[0][65] = 16'sd17;
        fc2_weights[0][66] = 16'sd3;
        fc2_weights[0][67] = 16'sd-49;
        fc2_weights[0][68] = 16'sd0;
        fc2_weights[0][69] = 16'sd106;
        fc2_weights[0][70] = 16'sd-67;
        fc2_weights[0][71] = 16'sd-11;
        fc2_weights[0][72] = 16'sd-31;
        fc2_weights[0][73] = 16'sd-51;
        fc2_weights[0][74] = 16'sd36;
        fc2_weights[0][75] = 16'sd19;
        fc2_weights[0][76] = 16'sd16;
        fc2_weights[0][77] = 16'sd-7;
        fc2_weights[0][78] = 16'sd4;
        fc2_weights[0][79] = 16'sd2;
        fc2_weights[0][80] = 16'sd-94;
        fc2_weights[0][81] = 16'sd-36;
        fc2_weights[0][82] = 16'sd-31;
        fc2_weights[0][83] = 16'sd-51;
        fc2_weights[0][84] = 16'sd69;
        fc2_weights[0][85] = 16'sd9;
        fc2_weights[0][86] = 16'sd-38;
        fc2_weights[0][87] = 16'sd-20;
        fc2_weights[0][88] = 16'sd46;
        fc2_weights[0][89] = 16'sd-78;
        fc2_weights[0][90] = 16'sd54;
        fc2_weights[0][91] = 16'sd-15;
        fc2_weights[0][92] = 16'sd18;
        fc2_weights[0][93] = 16'sd-17;
        fc2_weights[0][94] = 16'sd4;
        fc2_weights[0][95] = 16'sd-37;
        fc2_weights[0][96] = 16'sd97;
        fc2_weights[0][97] = 16'sd-20;
        fc2_weights[0][98] = 16'sd14;
        fc2_weights[0][99] = 16'sd-30;
        fc2_weights[0][100] = 16'sd37;
        fc2_weights[0][101] = 16'sd-28;
        fc2_weights[0][102] = 16'sd-2;
        fc2_weights[0][103] = 16'sd24;
        fc2_weights[0][104] = 16'sd31;
        fc2_weights[0][105] = 16'sd-34;
        fc2_weights[0][106] = 16'sd-2;
        fc2_weights[0][107] = 16'sd71;
        fc2_weights[0][108] = 16'sd-66;
        fc2_weights[0][109] = 16'sd10;
        fc2_weights[0][110] = 16'sd42;
        fc2_weights[0][111] = 16'sd-10;
        fc2_weights[0][112] = 16'sd1;
        fc2_weights[0][113] = 16'sd-72;
        fc2_weights[0][114] = 16'sd23;
        fc2_weights[0][115] = 16'sd-41;
        fc2_weights[0][116] = 16'sd9;
        fc2_weights[0][117] = 16'sd11;
        fc2_weights[0][118] = 16'sd-56;
        fc2_weights[0][119] = 16'sd9;
        fc2_weights[0][120] = 16'sd-57;
        fc2_weights[0][121] = 16'sd-20;
        fc2_weights[0][122] = 16'sd10;
        fc2_weights[0][123] = 16'sd39;
        fc2_weights[0][124] = 16'sd7;
        fc2_weights[0][125] = 16'sd64;
        fc2_weights[0][126] = 16'sd29;
        fc2_weights[0][127] = 16'sd-60;
        fc2_weights[1][0] = 16'sd-69;
        fc2_weights[1][1] = 16'sd-18;
        fc2_weights[1][2] = 16'sd-13;
        fc2_weights[1][3] = 16'sd-53;
        fc2_weights[1][4] = 16'sd47;
        fc2_weights[1][5] = 16'sd-15;
        fc2_weights[1][6] = 16'sd-14;
        fc2_weights[1][7] = 16'sd16;
        fc2_weights[1][8] = 16'sd27;
        fc2_weights[1][9] = 16'sd-37;
        fc2_weights[1][10] = 16'sd5;
        fc2_weights[1][11] = 16'sd32;
        fc2_weights[1][12] = 16'sd-13;
        fc2_weights[1][13] = 16'sd-19;
        fc2_weights[1][14] = 16'sd2;
        fc2_weights[1][15] = 16'sd-45;
        fc2_weights[1][16] = 16'sd44;
        fc2_weights[1][17] = 16'sd-23;
        fc2_weights[1][18] = 16'sd-84;
        fc2_weights[1][19] = 16'sd-8;
        fc2_weights[1][20] = 16'sd-85;
        fc2_weights[1][21] = 16'sd-31;
        fc2_weights[1][22] = 16'sd59;
        fc2_weights[1][23] = 16'sd38;
        fc2_weights[1][24] = 16'sd8;
        fc2_weights[1][25] = 16'sd-10;
        fc2_weights[1][26] = 16'sd8;
        fc2_weights[1][27] = 16'sd-19;
        fc2_weights[1][28] = 16'sd-26;
        fc2_weights[1][29] = 16'sd19;
        fc2_weights[1][30] = 16'sd-7;
        fc2_weights[1][31] = 16'sd-5;
        fc2_weights[1][32] = 16'sd-69;
        fc2_weights[1][33] = 16'sd-39;
        fc2_weights[1][34] = 16'sd-31;
        fc2_weights[1][35] = 16'sd-67;
        fc2_weights[1][36] = 16'sd79;
        fc2_weights[1][37] = 16'sd-61;
        fc2_weights[1][38] = 16'sd92;
        fc2_weights[1][39] = 16'sd19;
        fc2_weights[1][40] = 16'sd-94;
        fc2_weights[1][41] = 16'sd107;
        fc2_weights[1][42] = 16'sd38;
        fc2_weights[1][43] = 16'sd-45;
        fc2_weights[1][44] = 16'sd-9;
        fc2_weights[1][45] = 16'sd66;
        fc2_weights[1][46] = 16'sd20;
        fc2_weights[1][47] = 16'sd29;
        fc2_weights[1][48] = 16'sd19;
        fc2_weights[1][49] = 16'sd71;
        fc2_weights[1][50] = 16'sd-44;
        fc2_weights[1][51] = 16'sd79;
        fc2_weights[1][52] = 16'sd9;
        fc2_weights[1][53] = 16'sd38;
        fc2_weights[1][54] = 16'sd43;
        fc2_weights[1][55] = 16'sd12;
        fc2_weights[1][56] = 16'sd25;
        fc2_weights[1][57] = 16'sd-23;
        fc2_weights[1][58] = 16'sd-24;
        fc2_weights[1][59] = 16'sd-36;
        fc2_weights[1][60] = 16'sd38;
        fc2_weights[1][61] = 16'sd-47;
        fc2_weights[1][62] = 16'sd85;
        fc2_weights[1][63] = 16'sd-21;
        fc2_weights[1][64] = 16'sd70;
        fc2_weights[1][65] = 16'sd-8;
        fc2_weights[1][66] = 16'sd36;
        fc2_weights[1][67] = 16'sd0;
        fc2_weights[1][68] = 16'sd-18;
        fc2_weights[1][69] = 16'sd-61;
        fc2_weights[1][70] = 16'sd126;
        fc2_weights[1][71] = 16'sd-20;
        fc2_weights[1][72] = 16'sd-63;
        fc2_weights[1][73] = 16'sd11;
        fc2_weights[1][74] = 16'sd0;
        fc2_weights[1][75] = 16'sd-6;
        fc2_weights[1][76] = 16'sd19;
        fc2_weights[1][77] = 16'sd94;
        fc2_weights[1][78] = 16'sd-19;
        fc2_weights[1][79] = 16'sd29;
        fc2_weights[1][80] = 16'sd-52;
        fc2_weights[1][81] = 16'sd-8;
        fc2_weights[1][82] = 16'sd22;
        fc2_weights[1][83] = 16'sd-12;
        fc2_weights[1][84] = 16'sd-68;
        fc2_weights[1][85] = 16'sd3;
        fc2_weights[1][86] = 16'sd35;
        fc2_weights[1][87] = 16'sd-12;
        fc2_weights[1][88] = 16'sd39;
        fc2_weights[1][89] = 16'sd54;
        fc2_weights[1][90] = 16'sd-10;
        fc2_weights[1][91] = 16'sd55;
        fc2_weights[1][92] = 16'sd45;
        fc2_weights[1][93] = 16'sd24;
        fc2_weights[1][94] = 16'sd-109;
        fc2_weights[1][95] = 16'sd22;
        fc2_weights[1][96] = 16'sd-14;
        fc2_weights[1][97] = 16'sd-1;
        fc2_weights[1][98] = 16'sd2;
        fc2_weights[1][99] = 16'sd16;
        fc2_weights[1][100] = 16'sd-4;
        fc2_weights[1][101] = 16'sd7;
        fc2_weights[1][102] = 16'sd1;
        fc2_weights[1][103] = 16'sd-31;
        fc2_weights[1][104] = 16'sd32;
        fc2_weights[1][105] = 16'sd-61;
        fc2_weights[1][106] = 16'sd-14;
        fc2_weights[1][107] = 16'sd64;
        fc2_weights[1][108] = 16'sd0;
        fc2_weights[1][109] = 16'sd48;
        fc2_weights[1][110] = 16'sd3;
        fc2_weights[1][111] = 16'sd42;
        fc2_weights[1][112] = 16'sd-65;
        fc2_weights[1][113] = 16'sd16;
        fc2_weights[1][114] = 16'sd-16;
        fc2_weights[1][115] = 16'sd31;
        fc2_weights[1][116] = 16'sd-22;
        fc2_weights[1][117] = 16'sd-94;
        fc2_weights[1][118] = 16'sd76;
        fc2_weights[1][119] = 16'sd-26;
        fc2_weights[1][120] = 16'sd-28;
        fc2_weights[1][121] = 16'sd46;
        fc2_weights[1][122] = 16'sd11;
        fc2_weights[1][123] = 16'sd24;
        fc2_weights[1][124] = 16'sd-6;
        fc2_weights[1][125] = 16'sd-38;
        fc2_weights[1][126] = 16'sd34;
        fc2_weights[1][127] = 16'sd-43;
        fc2_weights[2][0] = 16'sd-51;
        fc2_weights[2][1] = 16'sd22;
        fc2_weights[2][2] = 16'sd31;
        fc2_weights[2][3] = 16'sd-36;
        fc2_weights[2][4] = 16'sd-14;
        fc2_weights[2][5] = 16'sd-7;
        fc2_weights[2][6] = 16'sd44;
        fc2_weights[2][7] = 16'sd-30;
        fc2_weights[2][8] = 16'sd35;
        fc2_weights[2][9] = 16'sd14;
        fc2_weights[2][10] = 16'sd-11;
        fc2_weights[2][11] = 16'sd-8;
        fc2_weights[2][12] = 16'sd-7;
        fc2_weights[2][13] = 16'sd-24;
        fc2_weights[2][14] = 16'sd-28;
        fc2_weights[2][15] = 16'sd5;
        fc2_weights[2][16] = 16'sd-35;
        fc2_weights[2][17] = 16'sd7;
        fc2_weights[2][18] = 16'sd-39;
        fc2_weights[2][19] = 16'sd-15;
        fc2_weights[2][20] = 16'sd3;
        fc2_weights[2][21] = 16'sd-24;
        fc2_weights[2][22] = 16'sd-30;
        fc2_weights[2][23] = 16'sd-25;
        fc2_weights[2][24] = 16'sd7;
        fc2_weights[2][25] = 16'sd27;
        fc2_weights[2][26] = 16'sd-6;
        fc2_weights[2][27] = 16'sd12;
        fc2_weights[2][28] = 16'sd-30;
        fc2_weights[2][29] = 16'sd-5;
        fc2_weights[2][30] = 16'sd10;
        fc2_weights[2][31] = 16'sd43;
        fc2_weights[2][32] = 16'sd0;
        fc2_weights[2][33] = 16'sd4;
        fc2_weights[2][34] = 16'sd35;
        fc2_weights[2][35] = 16'sd7;
        fc2_weights[2][36] = 16'sd-18;
        fc2_weights[2][37] = 16'sd-20;
        fc2_weights[2][38] = 16'sd72;
        fc2_weights[2][39] = 16'sd-21;
        fc2_weights[2][40] = 16'sd-45;
        fc2_weights[2][41] = 16'sd127;
        fc2_weights[2][42] = 16'sd-11;
        fc2_weights[2][43] = 16'sd-21;
        fc2_weights[2][44] = 16'sd-27;
        fc2_weights[2][45] = 16'sd17;
        fc2_weights[2][46] = 16'sd-32;
        fc2_weights[2][47] = 16'sd23;
        fc2_weights[2][48] = 16'sd39;
        fc2_weights[2][49] = 16'sd-8;
        fc2_weights[2][50] = 16'sd47;
        fc2_weights[2][51] = 16'sd18;
        fc2_weights[2][52] = 16'sd-14;
        fc2_weights[2][53] = 16'sd13;
        fc2_weights[2][54] = 16'sd57;
        fc2_weights[2][55] = 16'sd2;
        fc2_weights[2][56] = 16'sd-42;
        fc2_weights[2][57] = 16'sd-36;
        fc2_weights[2][58] = 16'sd20;
        fc2_weights[2][59] = 16'sd-10;
        fc2_weights[2][60] = 16'sd-28;
        fc2_weights[2][61] = 16'sd-35;
        fc2_weights[2][62] = 16'sd-34;
        fc2_weights[2][63] = 16'sd22;
        fc2_weights[2][64] = 16'sd2;
        fc2_weights[2][65] = 16'sd-88;
        fc2_weights[2][66] = 16'sd-27;
        fc2_weights[2][67] = 16'sd-15;
        fc2_weights[2][68] = 16'sd-15;
        fc2_weights[2][69] = 16'sd-23;
        fc2_weights[2][70] = 16'sd52;
        fc2_weights[2][71] = 16'sd-15;
        fc2_weights[2][72] = 16'sd29;
        fc2_weights[2][73] = 16'sd-37;
        fc2_weights[2][74] = 16'sd-18;
        fc2_weights[2][75] = 16'sd22;
        fc2_weights[2][76] = 16'sd15;
        fc2_weights[2][77] = 16'sd3;
        fc2_weights[2][78] = 16'sd5;
        fc2_weights[2][79] = 16'sd-29;
        fc2_weights[2][80] = 16'sd29;
        fc2_weights[2][81] = 16'sd-10;
        fc2_weights[2][82] = 16'sd-21;
        fc2_weights[2][83] = 16'sd12;
        fc2_weights[2][84] = 16'sd26;
        fc2_weights[2][85] = 16'sd-3;
        fc2_weights[2][86] = 16'sd16;
        fc2_weights[2][87] = 16'sd-45;
        fc2_weights[2][88] = 16'sd23;
        fc2_weights[2][89] = 16'sd-21;
        fc2_weights[2][90] = 16'sd0;
        fc2_weights[2][91] = 16'sd-11;
        fc2_weights[2][92] = 16'sd57;
        fc2_weights[2][93] = 16'sd-20;
        fc2_weights[2][94] = 16'sd-37;
        fc2_weights[2][95] = 16'sd26;
        fc2_weights[2][96] = 16'sd-21;
        fc2_weights[2][97] = 16'sd103;
        fc2_weights[2][98] = 16'sd-16;
        fc2_weights[2][99] = 16'sd18;
        fc2_weights[2][100] = 16'sd18;
        fc2_weights[2][101] = 16'sd-38;
        fc2_weights[2][102] = 16'sd-1;
        fc2_weights[2][103] = 16'sd7;
        fc2_weights[2][104] = 16'sd-36;
        fc2_weights[2][105] = 16'sd13;
        fc2_weights[2][106] = 16'sd35;
        fc2_weights[2][107] = 16'sd58;
        fc2_weights[2][108] = 16'sd-44;
        fc2_weights[2][109] = 16'sd-10;
        fc2_weights[2][110] = 16'sd50;
        fc2_weights[2][111] = 16'sd-15;
        fc2_weights[2][112] = 16'sd4;
        fc2_weights[2][113] = 16'sd-25;
        fc2_weights[2][114] = 16'sd-24;
        fc2_weights[2][115] = 16'sd-16;
        fc2_weights[2][116] = 16'sd33;
        fc2_weights[2][117] = 16'sd-32;
        fc2_weights[2][118] = 16'sd4;
        fc2_weights[2][119] = 16'sd15;
        fc2_weights[2][120] = 16'sd8;
        fc2_weights[2][121] = 16'sd138;
        fc2_weights[2][122] = 16'sd17;
        fc2_weights[2][123] = 16'sd-33;
        fc2_weights[2][124] = 16'sd59;
        fc2_weights[2][125] = 16'sd-10;
        fc2_weights[2][126] = 16'sd-11;
        fc2_weights[2][127] = 16'sd-45;
        fc2_weights[3][0] = 16'sd0;
        fc2_weights[3][1] = 16'sd8;
        fc2_weights[3][2] = 16'sd0;
        fc2_weights[3][3] = 16'sd61;
        fc2_weights[3][4] = 16'sd-97;
        fc2_weights[3][5] = 16'sd22;
        fc2_weights[3][6] = 16'sd-68;
        fc2_weights[3][7] = 16'sd-21;
        fc2_weights[3][8] = 16'sd-39;
        fc2_weights[3][9] = 16'sd11;
        fc2_weights[3][10] = 16'sd-15;
        fc2_weights[3][11] = 16'sd-75;
        fc2_weights[3][12] = 16'sd21;
        fc2_weights[3][13] = 16'sd6;
        fc2_weights[3][14] = 16'sd61;
        fc2_weights[3][15] = 16'sd43;
        fc2_weights[3][16] = 16'sd-24;
        fc2_weights[3][17] = 16'sd51;
        fc2_weights[3][18] = 16'sd-3;
        fc2_weights[3][19] = 16'sd-23;
        fc2_weights[3][20] = 16'sd28;
        fc2_weights[3][21] = 16'sd-21;
        fc2_weights[3][22] = 16'sd-15;
        fc2_weights[3][23] = 16'sd-18;
        fc2_weights[3][24] = 16'sd77;
        fc2_weights[3][25] = 16'sd-13;
        fc2_weights[3][26] = 16'sd4;
        fc2_weights[3][27] = 16'sd15;
        fc2_weights[3][28] = 16'sd1;
        fc2_weights[3][29] = 16'sd23;
        fc2_weights[3][30] = 16'sd-16;
        fc2_weights[3][31] = 16'sd-68;
        fc2_weights[3][32] = 16'sd60;
        fc2_weights[3][33] = 16'sd-58;
        fc2_weights[3][34] = 16'sd47;
        fc2_weights[3][35] = 16'sd20;
        fc2_weights[3][36] = 16'sd-66;
        fc2_weights[3][37] = 16'sd15;
        fc2_weights[3][38] = 16'sd-2;
        fc2_weights[3][39] = 16'sd-65;
        fc2_weights[3][40] = 16'sd47;
        fc2_weights[3][41] = 16'sd11;
        fc2_weights[3][42] = 16'sd-19;
        fc2_weights[3][43] = 16'sd-35;
        fc2_weights[3][44] = 16'sd59;
        fc2_weights[3][45] = 16'sd60;
        fc2_weights[3][46] = 16'sd-47;
        fc2_weights[3][47] = 16'sd12;
        fc2_weights[3][48] = 16'sd-7;
        fc2_weights[3][49] = 16'sd-2;
        fc2_weights[3][50] = 16'sd41;
        fc2_weights[3][51] = 16'sd-31;
        fc2_weights[3][52] = 16'sd30;
        fc2_weights[3][53] = 16'sd-58;
        fc2_weights[3][54] = 16'sd-102;
        fc2_weights[3][55] = 16'sd-1;
        fc2_weights[3][56] = 16'sd-19;
        fc2_weights[3][57] = 16'sd10;
        fc2_weights[3][58] = 16'sd3;
        fc2_weights[3][59] = 16'sd32;
        fc2_weights[3][60] = 16'sd48;
        fc2_weights[3][61] = 16'sd1;
        fc2_weights[3][62] = 16'sd19;
        fc2_weights[3][63] = 16'sd53;
        fc2_weights[3][64] = 16'sd-71;
        fc2_weights[3][65] = 16'sd60;
        fc2_weights[3][66] = 16'sd45;
        fc2_weights[3][67] = 16'sd-20;
        fc2_weights[3][68] = 16'sd16;
        fc2_weights[3][69] = 16'sd109;
        fc2_weights[3][70] = 16'sd19;
        fc2_weights[3][71] = 16'sd37;
        fc2_weights[3][72] = 16'sd-24;
        fc2_weights[3][73] = 16'sd-27;
        fc2_weights[3][74] = 16'sd57;
        fc2_weights[3][75] = 16'sd-32;
        fc2_weights[3][76] = 16'sd27;
        fc2_weights[3][77] = 16'sd-24;
        fc2_weights[3][78] = 16'sd-54;
        fc2_weights[3][79] = 16'sd-1;
        fc2_weights[3][80] = 16'sd-32;
        fc2_weights[3][81] = 16'sd-16;
        fc2_weights[3][82] = 16'sd-27;
        fc2_weights[3][83] = 16'sd-30;
        fc2_weights[3][84] = 16'sd59;
        fc2_weights[3][85] = 16'sd-30;
        fc2_weights[3][86] = 16'sd25;
        fc2_weights[3][87] = 16'sd-27;
        fc2_weights[3][88] = 16'sd27;
        fc2_weights[3][89] = 16'sd19;
        fc2_weights[3][90] = 16'sd79;
        fc2_weights[3][91] = 16'sd-14;
        fc2_weights[3][92] = 16'sd28;
        fc2_weights[3][93] = 16'sd-12;
        fc2_weights[3][94] = 16'sd35;
        fc2_weights[3][95] = 16'sd-4;
        fc2_weights[3][96] = 16'sd57;
        fc2_weights[3][97] = 16'sd-36;
        fc2_weights[3][98] = 16'sd-28;
        fc2_weights[3][99] = 16'sd-27;
        fc2_weights[3][100] = 16'sd5;
        fc2_weights[3][101] = 16'sd43;
        fc2_weights[3][102] = 16'sd-13;
        fc2_weights[3][103] = 16'sd-67;
        fc2_weights[3][104] = 16'sd2;
        fc2_weights[3][105] = 16'sd1;
        fc2_weights[3][106] = 16'sd-70;
        fc2_weights[3][107] = 16'sd1;
        fc2_weights[3][108] = 16'sd-39;
        fc2_weights[3][109] = 16'sd-6;
        fc2_weights[3][110] = 16'sd59;
        fc2_weights[3][111] = 16'sd-30;
        fc2_weights[3][112] = 16'sd0;
        fc2_weights[3][113] = 16'sd-95;
        fc2_weights[3][114] = 16'sd-1;
        fc2_weights[3][115] = 16'sd-68;
        fc2_weights[3][116] = 16'sd63;
        fc2_weights[3][117] = 16'sd67;
        fc2_weights[3][118] = 16'sd-70;
        fc2_weights[3][119] = 16'sd6;
        fc2_weights[3][120] = 16'sd-73;
        fc2_weights[3][121] = 16'sd-81;
        fc2_weights[3][122] = 16'sd60;
        fc2_weights[3][123] = 16'sd27;
        fc2_weights[3][124] = 16'sd-2;
        fc2_weights[3][125] = 16'sd34;
        fc2_weights[3][126] = 16'sd1;
        fc2_weights[3][127] = 16'sd43;
        fc2_weights[4][0] = 16'sd17;
        fc2_weights[4][1] = 16'sd-37;
        fc2_weights[4][2] = 16'sd16;
        fc2_weights[4][3] = 16'sd50;
        fc2_weights[4][4] = 16'sd-8;
        fc2_weights[4][5] = 16'sd-56;
        fc2_weights[4][6] = 16'sd-26;
        fc2_weights[4][7] = 16'sd8;
        fc2_weights[4][8] = 16'sd-30;
        fc2_weights[4][9] = 16'sd6;
        fc2_weights[4][10] = 16'sd-29;
        fc2_weights[4][11] = 16'sd-97;
        fc2_weights[4][12] = 16'sd12;
        fc2_weights[4][13] = 16'sd16;
        fc2_weights[4][14] = 16'sd26;
        fc2_weights[4][15] = 16'sd38;
        fc2_weights[4][16] = 16'sd48;
        fc2_weights[4][17] = 16'sd-3;
        fc2_weights[4][18] = 16'sd-45;
        fc2_weights[4][19] = 16'sd19;
        fc2_weights[4][20] = 16'sd-8;
        fc2_weights[4][21] = 16'sd-40;
        fc2_weights[4][22] = 16'sd-18;
        fc2_weights[4][23] = 16'sd-6;
        fc2_weights[4][24] = 16'sd-25;
        fc2_weights[4][25] = 16'sd-25;
        fc2_weights[4][26] = 16'sd6;
        fc2_weights[4][27] = 16'sd9;
        fc2_weights[4][28] = 16'sd19;
        fc2_weights[4][29] = 16'sd-8;
        fc2_weights[4][30] = 16'sd22;
        fc2_weights[4][31] = 16'sd-34;
        fc2_weights[4][32] = 16'sd-77;
        fc2_weights[4][33] = 16'sd-38;
        fc2_weights[4][34] = 16'sd44;
        fc2_weights[4][35] = 16'sd86;
        fc2_weights[4][36] = 16'sd-48;
        fc2_weights[4][37] = 16'sd32;
        fc2_weights[4][38] = 16'sd-13;
        fc2_weights[4][39] = 16'sd14;
        fc2_weights[4][40] = 16'sd38;
        fc2_weights[4][41] = 16'sd-3;
        fc2_weights[4][42] = 16'sd5;
        fc2_weights[4][43] = 16'sd-8;
        fc2_weights[4][44] = 16'sd35;
        fc2_weights[4][45] = 16'sd56;
        fc2_weights[4][46] = 16'sd-15;
        fc2_weights[4][47] = 16'sd-20;
        fc2_weights[4][48] = 16'sd26;
        fc2_weights[4][49] = 16'sd37;
        fc2_weights[4][50] = 16'sd-13;
        fc2_weights[4][51] = 16'sd2;
        fc2_weights[4][52] = 16'sd44;
        fc2_weights[4][53] = 16'sd-49;
        fc2_weights[4][54] = 16'sd13;
        fc2_weights[4][55] = 16'sd-25;
        fc2_weights[4][56] = 16'sd58;
        fc2_weights[4][57] = 16'sd75;
        fc2_weights[4][58] = 16'sd-4;
        fc2_weights[4][59] = 16'sd3;
        fc2_weights[4][60] = 16'sd0;
        fc2_weights[4][61] = 16'sd-10;
        fc2_weights[4][62] = 16'sd6;
        fc2_weights[4][63] = 16'sd-37;
        fc2_weights[4][64] = 16'sd-4;
        fc2_weights[4][65] = 16'sd2;
        fc2_weights[4][66] = 16'sd-8;
        fc2_weights[4][67] = 16'sd-88;
        fc2_weights[4][68] = 16'sd-9;
        fc2_weights[4][69] = 16'sd10;
        fc2_weights[4][70] = 16'sd9;
        fc2_weights[4][71] = 16'sd54;
        fc2_weights[4][72] = 16'sd-46;
        fc2_weights[4][73] = 16'sd-43;
        fc2_weights[4][74] = 16'sd-3;
        fc2_weights[4][75] = 16'sd16;
        fc2_weights[4][76] = 16'sd-12;
        fc2_weights[4][77] = 16'sd17;
        fc2_weights[4][78] = 16'sd13;
        fc2_weights[4][79] = 16'sd-40;
        fc2_weights[4][80] = 16'sd-22;
        fc2_weights[4][81] = 16'sd35;
        fc2_weights[4][82] = 16'sd-40;
        fc2_weights[4][83] = 16'sd5;
        fc2_weights[4][84] = 16'sd-57;
        fc2_weights[4][85] = 16'sd4;
        fc2_weights[4][86] = 16'sd20;
        fc2_weights[4][87] = 16'sd1;
        fc2_weights[4][88] = 16'sd22;
        fc2_weights[4][89] = 16'sd-36;
        fc2_weights[4][90] = 16'sd-14;
        fc2_weights[4][91] = 16'sd17;
        fc2_weights[4][92] = 16'sd-5;
        fc2_weights[4][93] = 16'sd-14;
        fc2_weights[4][94] = 16'sd11;
        fc2_weights[4][95] = 16'sd-34;
        fc2_weights[4][96] = 16'sd12;
        fc2_weights[4][97] = 16'sd-21;
        fc2_weights[4][98] = 16'sd34;
        fc2_weights[4][99] = 16'sd-30;
        fc2_weights[4][100] = 16'sd11;
        fc2_weights[4][101] = 16'sd21;
        fc2_weights[4][102] = 16'sd-8;
        fc2_weights[4][103] = 16'sd-2;
        fc2_weights[4][104] = 16'sd63;
        fc2_weights[4][105] = 16'sd-27;
        fc2_weights[4][106] = 16'sd-8;
        fc2_weights[4][107] = 16'sd-12;
        fc2_weights[4][108] = 16'sd-73;
        fc2_weights[4][109] = 16'sd-26;
        fc2_weights[4][110] = 16'sd35;
        fc2_weights[4][111] = 16'sd-12;
        fc2_weights[4][112] = 16'sd19;
        fc2_weights[4][113] = 16'sd-62;
        fc2_weights[4][114] = 16'sd-3;
        fc2_weights[4][115] = 16'sd-41;
        fc2_weights[4][116] = 16'sd1;
        fc2_weights[4][117] = 16'sd-25;
        fc2_weights[4][118] = 16'sd-40;
        fc2_weights[4][119] = 16'sd-18;
        fc2_weights[4][120] = 16'sd-38;
        fc2_weights[4][121] = 16'sd-61;
        fc2_weights[4][122] = 16'sd-39;
        fc2_weights[4][123] = 16'sd27;
        fc2_weights[4][124] = 16'sd-54;
        fc2_weights[4][125] = 16'sd11;
        fc2_weights[4][126] = 16'sd-4;
        fc2_weights[4][127] = 16'sd-3;
        fc2_weights[5][0] = 16'sd-14;
        fc2_weights[5][1] = 16'sd-38;
        fc2_weights[5][2] = 16'sd-19;
        fc2_weights[5][3] = 16'sd25;
        fc2_weights[5][4] = 16'sd-16;
        fc2_weights[5][5] = 16'sd12;
        fc2_weights[5][6] = 16'sd-18;
        fc2_weights[5][7] = 16'sd4;
        fc2_weights[5][8] = 16'sd-10;
        fc2_weights[5][9] = 16'sd2;
        fc2_weights[5][10] = 16'sd31;
        fc2_weights[5][11] = 16'sd1;
        fc2_weights[5][12] = 16'sd-1;
        fc2_weights[5][13] = 16'sd46;
        fc2_weights[5][14] = 16'sd-13;
        fc2_weights[5][15] = 16'sd-1;
        fc2_weights[5][16] = 16'sd-14;
        fc2_weights[5][17] = 16'sd30;
        fc2_weights[5][18] = 16'sd-6;
        fc2_weights[5][19] = 16'sd30;
        fc2_weights[5][20] = 16'sd10;
        fc2_weights[5][21] = 16'sd11;
        fc2_weights[5][22] = 16'sd5;
        fc2_weights[5][23] = 16'sd5;
        fc2_weights[5][24] = 16'sd30;
        fc2_weights[5][25] = 16'sd2;
        fc2_weights[5][26] = 16'sd-1;
        fc2_weights[5][27] = 16'sd11;
        fc2_weights[5][28] = 16'sd-5;
        fc2_weights[5][29] = 16'sd7;
        fc2_weights[5][30] = 16'sd30;
        fc2_weights[5][31] = 16'sd-34;
        fc2_weights[5][32] = 16'sd4;
        fc2_weights[5][33] = 16'sd-24;
        fc2_weights[5][34] = 16'sd23;
        fc2_weights[5][35] = 16'sd4;
        fc2_weights[5][36] = 16'sd-1;
        fc2_weights[5][37] = 16'sd-1;
        fc2_weights[5][38] = 16'sd-27;
        fc2_weights[5][39] = 16'sd-21;
        fc2_weights[5][40] = 16'sd21;
        fc2_weights[5][41] = 16'sd-17;
        fc2_weights[5][42] = 16'sd12;
        fc2_weights[5][43] = 16'sd14;
        fc2_weights[5][44] = 16'sd12;
        fc2_weights[5][45] = 16'sd27;
        fc2_weights[5][46] = 16'sd-28;
        fc2_weights[5][47] = 16'sd-23;
        fc2_weights[5][48] = 16'sd41;
        fc2_weights[5][49] = 16'sd-2;
        fc2_weights[5][50] = 16'sd21;
        fc2_weights[5][51] = 16'sd40;
        fc2_weights[5][52] = 16'sd44;
        fc2_weights[5][53] = 16'sd14;
        fc2_weights[5][54] = 16'sd-27;
        fc2_weights[5][55] = 16'sd-13;
        fc2_weights[5][56] = 16'sd26;
        fc2_weights[5][57] = 16'sd23;
        fc2_weights[5][58] = 16'sd20;
        fc2_weights[5][59] = 16'sd39;
        fc2_weights[5][60] = 16'sd13;
        fc2_weights[5][61] = 16'sd22;
        fc2_weights[5][62] = 16'sd1;
        fc2_weights[5][63] = 16'sd21;
        fc2_weights[5][64] = 16'sd-25;
        fc2_weights[5][65] = 16'sd31;
        fc2_weights[5][66] = 16'sd33;
        fc2_weights[5][67] = 16'sd-43;
        fc2_weights[5][68] = 16'sd-11;
        fc2_weights[5][69] = 16'sd8;
        fc2_weights[5][70] = 16'sd-23;
        fc2_weights[5][71] = 16'sd21;
        fc2_weights[5][72] = 16'sd-19;
        fc2_weights[5][73] = 16'sd-19;
        fc2_weights[5][74] = 16'sd2;
        fc2_weights[5][75] = 16'sd7;
        fc2_weights[5][76] = 16'sd-3;
        fc2_weights[5][77] = 16'sd-9;
        fc2_weights[5][78] = 16'sd23;
        fc2_weights[5][79] = 16'sd-17;
        fc2_weights[5][80] = 16'sd-50;
        fc2_weights[5][81] = 16'sd-15;
        fc2_weights[5][82] = 16'sd-32;
        fc2_weights[5][83] = 16'sd-6;
        fc2_weights[5][84] = 16'sd3;
        fc2_weights[5][85] = 16'sd16;
        fc2_weights[5][86] = 16'sd-23;
        fc2_weights[5][87] = 16'sd-24;
        fc2_weights[5][88] = 16'sd14;
        fc2_weights[5][89] = 16'sd-53;
        fc2_weights[5][90] = 16'sd26;
        fc2_weights[5][91] = 16'sd6;
        fc2_weights[5][92] = 16'sd18;
        fc2_weights[5][93] = 16'sd-4;
        fc2_weights[5][94] = 16'sd-16;
        fc2_weights[5][95] = 16'sd-15;
        fc2_weights[5][96] = 16'sd19;
        fc2_weights[5][97] = 16'sd-2;
        fc2_weights[5][98] = 16'sd-16;
        fc2_weights[5][99] = 16'sd-18;
        fc2_weights[5][100] = 16'sd16;
        fc2_weights[5][101] = 16'sd-11;
        fc2_weights[5][102] = 16'sd-8;
        fc2_weights[5][103] = 16'sd35;
        fc2_weights[5][104] = 16'sd3;
        fc2_weights[5][105] = 16'sd3;
        fc2_weights[5][106] = 16'sd-27;
        fc2_weights[5][107] = 16'sd1;
        fc2_weights[5][108] = 16'sd-35;
        fc2_weights[5][109] = 16'sd-25;
        fc2_weights[5][110] = 16'sd31;
        fc2_weights[5][111] = 16'sd-31;
        fc2_weights[5][112] = 16'sd-28;
        fc2_weights[5][113] = 16'sd-22;
        fc2_weights[5][114] = 16'sd-3;
        fc2_weights[5][115] = 16'sd10;
        fc2_weights[5][116] = 16'sd-1;
        fc2_weights[5][117] = 16'sd1;
        fc2_weights[5][118] = 16'sd-43;
        fc2_weights[5][119] = 16'sd6;
        fc2_weights[5][120] = 16'sd-24;
        fc2_weights[5][121] = 16'sd3;
        fc2_weights[5][122] = 16'sd19;
        fc2_weights[5][123] = 16'sd23;
        fc2_weights[5][124] = 16'sd-3;
        fc2_weights[5][125] = 16'sd36;
        fc2_weights[5][126] = 16'sd32;
        fc2_weights[5][127] = 16'sd60;
        fc2_weights[6][0] = 16'sd-2;
        fc2_weights[6][1] = 16'sd16;
        fc2_weights[6][2] = 16'sd-67;
        fc2_weights[6][3] = 16'sd2;
        fc2_weights[6][4] = 16'sd39;
        fc2_weights[6][5] = 16'sd1;
        fc2_weights[6][6] = 16'sd-21;
        fc2_weights[6][7] = 16'sd21;
        fc2_weights[6][8] = 16'sd50;
        fc2_weights[6][9] = 16'sd3;
        fc2_weights[6][10] = 16'sd-22;
        fc2_weights[6][11] = 16'sd29;
        fc2_weights[6][12] = 16'sd82;
        fc2_weights[6][13] = 16'sd-13;
        fc2_weights[6][14] = 16'sd-35;
        fc2_weights[6][15] = 16'sd-3;
        fc2_weights[6][16] = 16'sd-20;
        fc2_weights[6][17] = 16'sd3;
        fc2_weights[6][18] = 16'sd-4;
        fc2_weights[6][19] = 16'sd-40;
        fc2_weights[6][20] = 16'sd-21;
        fc2_weights[6][21] = 16'sd-18;
        fc2_weights[6][22] = 16'sd-4;
        fc2_weights[6][23] = 16'sd-8;
        fc2_weights[6][24] = 16'sd-8;
        fc2_weights[6][25] = 16'sd-62;
        fc2_weights[6][26] = 16'sd-5;
        fc2_weights[6][27] = 16'sd-21;
        fc2_weights[6][28] = 16'sd15;
        fc2_weights[6][29] = 16'sd-58;
        fc2_weights[6][30] = 16'sd-21;
        fc2_weights[6][31] = 16'sd72;
        fc2_weights[6][32] = 16'sd17;
        fc2_weights[6][33] = 16'sd59;
        fc2_weights[6][34] = 16'sd-24;
        fc2_weights[6][35] = 16'sd-22;
        fc2_weights[6][36] = 16'sd-4;
        fc2_weights[6][37] = 16'sd20;
        fc2_weights[6][38] = 16'sd-26;
        fc2_weights[6][39] = 16'sd36;
        fc2_weights[6][40] = 16'sd48;
        fc2_weights[6][41] = 16'sd-18;
        fc2_weights[6][42] = 16'sd-56;
        fc2_weights[6][43] = 16'sd11;
        fc2_weights[6][44] = 16'sd4;
        fc2_weights[6][45] = 16'sd-42;
        fc2_weights[6][46] = 16'sd-47;
        fc2_weights[6][47] = 16'sd-15;
        fc2_weights[6][48] = 16'sd-55;
        fc2_weights[6][49] = 16'sd7;
        fc2_weights[6][50] = 16'sd-13;
        fc2_weights[6][51] = 16'sd-79;
        fc2_weights[6][52] = 16'sd-40;
        fc2_weights[6][53] = 16'sd-36;
        fc2_weights[6][54] = 16'sd-8;
        fc2_weights[6][55] = 16'sd-12;
        fc2_weights[6][56] = 16'sd-17;
        fc2_weights[6][57] = 16'sd-24;
        fc2_weights[6][58] = 16'sd-31;
        fc2_weights[6][59] = 16'sd-32;
        fc2_weights[6][60] = 16'sd-44;
        fc2_weights[6][61] = 16'sd24;
        fc2_weights[6][62] = 16'sd-48;
        fc2_weights[6][63] = 16'sd-5;
        fc2_weights[6][64] = 16'sd-20;
        fc2_weights[6][65] = 16'sd-55;
        fc2_weights[6][66] = 16'sd-44;
        fc2_weights[6][67] = 16'sd17;
        fc2_weights[6][68] = 16'sd42;
        fc2_weights[6][69] = 16'sd9;
        fc2_weights[6][70] = 16'sd33;
        fc2_weights[6][71] = 16'sd-23;
        fc2_weights[6][72] = 16'sd5;
        fc2_weights[6][73] = 16'sd24;
        fc2_weights[6][74] = 16'sd-31;
        fc2_weights[6][75] = 16'sd-35;
        fc2_weights[6][76] = 16'sd-2;
        fc2_weights[6][77] = 16'sd2;
        fc2_weights[6][78] = 16'sd21;
        fc2_weights[6][79] = 16'sd-4;
        fc2_weights[6][80] = 16'sd-28;
        fc2_weights[6][81] = 16'sd-73;
        fc2_weights[6][82] = 16'sd-18;
        fc2_weights[6][83] = 16'sd31;
        fc2_weights[6][84] = 16'sd9;
        fc2_weights[6][85] = 16'sd-22;
        fc2_weights[6][86] = 16'sd-14;
        fc2_weights[6][87] = 16'sd38;
        fc2_weights[6][88] = 16'sd0;
        fc2_weights[6][89] = 16'sd25;
        fc2_weights[6][90] = 16'sd-38;
        fc2_weights[6][91] = 16'sd16;
        fc2_weights[6][92] = 16'sd-3;
        fc2_weights[6][93] = 16'sd48;
        fc2_weights[6][94] = 16'sd1;
        fc2_weights[6][95] = 16'sd-1;
        fc2_weights[6][96] = 16'sd-8;
        fc2_weights[6][97] = 16'sd-3;
        fc2_weights[6][98] = 16'sd-44;
        fc2_weights[6][99] = 16'sd14;
        fc2_weights[6][100] = 16'sd-30;
        fc2_weights[6][101] = 16'sd2;
        fc2_weights[6][102] = 16'sd-21;
        fc2_weights[6][103] = 16'sd-31;
        fc2_weights[6][104] = 16'sd-20;
        fc2_weights[6][105] = 16'sd-33;
        fc2_weights[6][106] = 16'sd-7;
        fc2_weights[6][107] = 16'sd-43;
        fc2_weights[6][108] = 16'sd-86;
        fc2_weights[6][109] = 16'sd-15;
        fc2_weights[6][110] = 16'sd-42;
        fc2_weights[6][111] = 16'sd-48;
        fc2_weights[6][112] = 16'sd30;
        fc2_weights[6][113] = 16'sd-6;
        fc2_weights[6][114] = 16'sd15;
        fc2_weights[6][115] = 16'sd-11;
        fc2_weights[6][116] = 16'sd-22;
        fc2_weights[6][117] = 16'sd7;
        fc2_weights[6][118] = 16'sd-23;
        fc2_weights[6][119] = 16'sd25;
        fc2_weights[6][120] = 16'sd31;
        fc2_weights[6][121] = 16'sd-24;
        fc2_weights[6][122] = 16'sd3;
        fc2_weights[6][123] = 16'sd-18;
        fc2_weights[6][124] = 16'sd9;
        fc2_weights[6][125] = 16'sd-49;
        fc2_weights[6][126] = 16'sd-37;
        fc2_weights[6][127] = 16'sd-87;
        fc2_weights[7][0] = 16'sd-3;
        fc2_weights[7][1] = 16'sd-52;
        fc2_weights[7][2] = 16'sd48;
        fc2_weights[7][3] = 16'sd-58;
        fc2_weights[7][4] = 16'sd-6;
        fc2_weights[7][5] = 16'sd-7;
        fc2_weights[7][6] = 16'sd54;
        fc2_weights[7][7] = 16'sd25;
        fc2_weights[7][8] = 16'sd39;
        fc2_weights[7][9] = 16'sd-28;
        fc2_weights[7][10] = 16'sd-38;
        fc2_weights[7][11] = 16'sd23;
        fc2_weights[7][12] = 16'sd-43;
        fc2_weights[7][13] = 16'sd-11;
        fc2_weights[7][14] = 16'sd55;
        fc2_weights[7][15] = 16'sd-50;
        fc2_weights[7][16] = 16'sd37;
        fc2_weights[7][17] = 16'sd-64;
        fc2_weights[7][18] = 16'sd0;
        fc2_weights[7][19] = 16'sd27;
        fc2_weights[7][20] = 16'sd22;
        fc2_weights[7][21] = 16'sd12;
        fc2_weights[7][22] = 16'sd-10;
        fc2_weights[7][23] = 16'sd20;
        fc2_weights[7][24] = 16'sd14;
        fc2_weights[7][25] = 16'sd4;
        fc2_weights[7][26] = 16'sd-20;
        fc2_weights[7][27] = 16'sd-10;
        fc2_weights[7][28] = 16'sd-5;
        fc2_weights[7][29] = 16'sd5;
        fc2_weights[7][30] = 16'sd-68;
        fc2_weights[7][31] = 16'sd3;
        fc2_weights[7][32] = 16'sd-54;
        fc2_weights[7][33] = 16'sd-27;
        fc2_weights[7][34] = 16'sd-33;
        fc2_weights[7][35] = 16'sd3;
        fc2_weights[7][36] = 16'sd-64;
        fc2_weights[7][37] = 16'sd-68;
        fc2_weights[7][38] = 16'sd16;
        fc2_weights[7][39] = 16'sd-7;
        fc2_weights[7][40] = 16'sd-7;
        fc2_weights[7][41] = 16'sd100;
        fc2_weights[7][42] = 16'sd-45;
        fc2_weights[7][43] = 16'sd10;
        fc2_weights[7][44] = 16'sd-11;
        fc2_weights[7][45] = 16'sd7;
        fc2_weights[7][46] = 16'sd57;
        fc2_weights[7][47] = 16'sd-22;
        fc2_weights[7][48] = 16'sd23;
        fc2_weights[7][49] = 16'sd52;
        fc2_weights[7][50] = 16'sd22;
        fc2_weights[7][51] = 16'sd-34;
        fc2_weights[7][52] = 16'sd22;
        fc2_weights[7][53] = 16'sd-54;
        fc2_weights[7][54] = 16'sd91;
        fc2_weights[7][55] = 16'sd53;
        fc2_weights[7][56] = 16'sd27;
        fc2_weights[7][57] = 16'sd-31;
        fc2_weights[7][58] = 16'sd-13;
        fc2_weights[7][59] = 16'sd5;
        fc2_weights[7][60] = 16'sd68;
        fc2_weights[7][61] = 16'sd-58;
        fc2_weights[7][62] = 16'sd8;
        fc2_weights[7][63] = 16'sd12;
        fc2_weights[7][64] = 16'sd40;
        fc2_weights[7][65] = 16'sd28;
        fc2_weights[7][66] = 16'sd15;
        fc2_weights[7][67] = 16'sd-8;
        fc2_weights[7][68] = 16'sd-14;
        fc2_weights[7][69] = 16'sd-55;
        fc2_weights[7][70] = 16'sd40;
        fc2_weights[7][71] = 16'sd51;
        fc2_weights[7][72] = 16'sd20;
        fc2_weights[7][73] = 16'sd23;
        fc2_weights[7][74] = 16'sd-2;
        fc2_weights[7][75] = 16'sd43;
        fc2_weights[7][76] = 16'sd-12;
        fc2_weights[7][77] = 16'sd31;
        fc2_weights[7][78] = 16'sd23;
        fc2_weights[7][79] = 16'sd49;
        fc2_weights[7][80] = 16'sd21;
        fc2_weights[7][81] = 16'sd18;
        fc2_weights[7][82] = 16'sd-31;
        fc2_weights[7][83] = 16'sd-25;
        fc2_weights[7][84] = 16'sd-64;
        fc2_weights[7][85] = 16'sd-14;
        fc2_weights[7][86] = 16'sd11;
        fc2_weights[7][87] = 16'sd-7;
        fc2_weights[7][88] = 16'sd40;
        fc2_weights[7][89] = 16'sd47;
        fc2_weights[7][90] = 16'sd1;
        fc2_weights[7][91] = 16'sd-13;
        fc2_weights[7][92] = 16'sd50;
        fc2_weights[7][93] = 16'sd-7;
        fc2_weights[7][94] = 16'sd-48;
        fc2_weights[7][95] = 16'sd-9;
        fc2_weights[7][96] = 16'sd-36;
        fc2_weights[7][97] = 16'sd54;
        fc2_weights[7][98] = 16'sd14;
        fc2_weights[7][99] = 16'sd19;
        fc2_weights[7][100] = 16'sd30;
        fc2_weights[7][101] = 16'sd-26;
        fc2_weights[7][102] = 16'sd55;
        fc2_weights[7][103] = 16'sd-13;
        fc2_weights[7][104] = 16'sd-11;
        fc2_weights[7][105] = 16'sd-8;
        fc2_weights[7][106] = 16'sd-24;
        fc2_weights[7][107] = 16'sd48;
        fc2_weights[7][108] = 16'sd-19;
        fc2_weights[7][109] = 16'sd6;
        fc2_weights[7][110] = 16'sd25;
        fc2_weights[7][111] = 16'sd39;
        fc2_weights[7][112] = 16'sd-41;
        fc2_weights[7][113] = 16'sd-16;
        fc2_weights[7][114] = 16'sd-16;
        fc2_weights[7][115] = 16'sd2;
        fc2_weights[7][116] = 16'sd-39;
        fc2_weights[7][117] = 16'sd-129;
        fc2_weights[7][118] = 16'sd-4;
        fc2_weights[7][119] = 16'sd-22;
        fc2_weights[7][120] = 16'sd21;
        fc2_weights[7][121] = 16'sd45;
        fc2_weights[7][122] = 16'sd1;
        fc2_weights[7][123] = 16'sd35;
        fc2_weights[7][124] = 16'sd43;
        fc2_weights[7][125] = 16'sd-22;
        fc2_weights[7][126] = 16'sd39;
        fc2_weights[7][127] = 16'sd-8;
        fc2_weights[8][0] = 16'sd23;
        fc2_weights[8][1] = 16'sd-23;
        fc2_weights[8][2] = 16'sd-13;
        fc2_weights[8][3] = 16'sd6;
        fc2_weights[8][4] = 16'sd8;
        fc2_weights[8][5] = 16'sd8;
        fc2_weights[8][6] = 16'sd-5;
        fc2_weights[8][7] = 16'sd34;
        fc2_weights[8][8] = 16'sd38;
        fc2_weights[8][9] = 16'sd29;
        fc2_weights[8][10] = 16'sd11;
        fc2_weights[8][11] = 16'sd6;
        fc2_weights[8][12] = 16'sd12;
        fc2_weights[8][13] = 16'sd-62;
        fc2_weights[8][14] = 16'sd-1;
        fc2_weights[8][15] = 16'sd-49;
        fc2_weights[8][16] = 16'sd30;
        fc2_weights[8][17] = 16'sd-102;
        fc2_weights[8][18] = 16'sd28;
        fc2_weights[8][19] = 16'sd-18;
        fc2_weights[8][20] = 16'sd-31;
        fc2_weights[8][21] = 16'sd-5;
        fc2_weights[8][22] = 16'sd37;
        fc2_weights[8][23] = 16'sd63;
        fc2_weights[8][24] = 16'sd-49;
        fc2_weights[8][25] = 16'sd-39;
        fc2_weights[8][26] = 16'sd20;
        fc2_weights[8][27] = 16'sd-6;
        fc2_weights[8][28] = 16'sd29;
        fc2_weights[8][29] = 16'sd20;
        fc2_weights[8][30] = 16'sd-51;
        fc2_weights[8][31] = 16'sd39;
        fc2_weights[8][32] = 16'sd-57;
        fc2_weights[8][33] = 16'sd-8;
        fc2_weights[8][34] = 16'sd-35;
        fc2_weights[8][35] = 16'sd15;
        fc2_weights[8][36] = 16'sd45;
        fc2_weights[8][37] = 16'sd29;
        fc2_weights[8][38] = 16'sd33;
        fc2_weights[8][39] = 16'sd32;
        fc2_weights[8][40] = 16'sd-23;
        fc2_weights[8][41] = 16'sd-37;
        fc2_weights[8][42] = 16'sd-21;
        fc2_weights[8][43] = 16'sd-2;
        fc2_weights[8][44] = 16'sd-21;
        fc2_weights[8][45] = 16'sd-4;
        fc2_weights[8][46] = 16'sd27;
        fc2_weights[8][47] = 16'sd-26;
        fc2_weights[8][48] = 16'sd-31;
        fc2_weights[8][49] = 16'sd-10;
        fc2_weights[8][50] = 16'sd-66;
        fc2_weights[8][51] = 16'sd40;
        fc2_weights[8][52] = 16'sd-63;
        fc2_weights[8][53] = 16'sd41;
        fc2_weights[8][54] = 16'sd53;
        fc2_weights[8][55] = 16'sd38;
        fc2_weights[8][56] = 16'sd-26;
        fc2_weights[8][57] = 16'sd-59;
        fc2_weights[8][58] = 16'sd-37;
        fc2_weights[8][59] = 16'sd-88;
        fc2_weights[8][60] = 16'sd35;
        fc2_weights[8][61] = 16'sd15;
        fc2_weights[8][62] = 16'sd11;
        fc2_weights[8][63] = 16'sd-62;
        fc2_weights[8][64] = 16'sd20;
        fc2_weights[8][65] = 16'sd-6;
        fc2_weights[8][66] = 16'sd-3;
        fc2_weights[8][67] = 16'sd22;
        fc2_weights[8][68] = 16'sd-5;
        fc2_weights[8][69] = 16'sd-74;
        fc2_weights[8][70] = 16'sd17;
        fc2_weights[8][71] = 16'sd-28;
        fc2_weights[8][72] = 16'sd20;
        fc2_weights[8][73] = 16'sd-21;
        fc2_weights[8][74] = 16'sd-13;
        fc2_weights[8][75] = 16'sd23;
        fc2_weights[8][76] = 16'sd34;
        fc2_weights[8][77] = 16'sd35;
        fc2_weights[8][78] = 16'sd-71;
        fc2_weights[8][79] = 16'sd-10;
        fc2_weights[8][80] = 16'sd-6;
        fc2_weights[8][81] = 16'sd11;
        fc2_weights[8][82] = 16'sd24;
        fc2_weights[8][83] = 16'sd43;
        fc2_weights[8][84] = 16'sd-31;
        fc2_weights[8][85] = 16'sd11;
        fc2_weights[8][86] = 16'sd-30;
        fc2_weights[8][87] = 16'sd-23;
        fc2_weights[8][88] = 16'sd-57;
        fc2_weights[8][89] = 16'sd42;
        fc2_weights[8][90] = 16'sd-54;
        fc2_weights[8][91] = 16'sd41;
        fc2_weights[8][92] = 16'sd25;
        fc2_weights[8][93] = 16'sd19;
        fc2_weights[8][94] = 16'sd-9;
        fc2_weights[8][95] = 16'sd38;
        fc2_weights[8][96] = 16'sd-69;
        fc2_weights[8][97] = 16'sd-16;
        fc2_weights[8][98] = 16'sd58;
        fc2_weights[8][99] = 16'sd34;
        fc2_weights[8][100] = 16'sd-46;
        fc2_weights[8][101] = 16'sd-22;
        fc2_weights[8][102] = 16'sd-4;
        fc2_weights[8][103] = 16'sd8;
        fc2_weights[8][104] = 16'sd11;
        fc2_weights[8][105] = 16'sd19;
        fc2_weights[8][106] = 16'sd-1;
        fc2_weights[8][107] = 16'sd10;
        fc2_weights[8][108] = 16'sd33;
        fc2_weights[8][109] = 16'sd1;
        fc2_weights[8][110] = 16'sd-61;
        fc2_weights[8][111] = 16'sd17;
        fc2_weights[8][112] = 16'sd-1;
        fc2_weights[8][113] = 16'sd-3;
        fc2_weights[8][114] = 16'sd-2;
        fc2_weights[8][115] = 16'sd49;
        fc2_weights[8][116] = 16'sd-22;
        fc2_weights[8][117] = 16'sd-100;
        fc2_weights[8][118] = 16'sd60;
        fc2_weights[8][119] = 16'sd-4;
        fc2_weights[8][120] = 16'sd16;
        fc2_weights[8][121] = 16'sd29;
        fc2_weights[8][122] = 16'sd-51;
        fc2_weights[8][123] = 16'sd-11;
        fc2_weights[8][124] = 16'sd-12;
        fc2_weights[8][125] = 16'sd-6;
        fc2_weights[8][126] = 16'sd-15;
        fc2_weights[8][127] = 16'sd-39;
        fc2_weights[9][0] = 16'sd-7;
        fc2_weights[9][1] = 16'sd-58;
        fc2_weights[9][2] = 16'sd10;
        fc2_weights[9][3] = 16'sd-30;
        fc2_weights[9][4] = 16'sd-2;
        fc2_weights[9][5] = 16'sd20;
        fc2_weights[9][6] = 16'sd-41;
        fc2_weights[9][7] = 16'sd-22;
        fc2_weights[9][8] = 16'sd-3;
        fc2_weights[9][9] = 16'sd-15;
        fc2_weights[9][10] = 16'sd7;
        fc2_weights[9][11] = 16'sd-54;
        fc2_weights[9][12] = 16'sd-21;
        fc2_weights[9][13] = 16'sd-23;
        fc2_weights[9][14] = 16'sd63;
        fc2_weights[9][15] = 16'sd25;
        fc2_weights[9][16] = 16'sd-25;
        fc2_weights[9][17] = 16'sd-30;
        fc2_weights[9][18] = 16'sd13;
        fc2_weights[9][19] = 16'sd16;
        fc2_weights[9][20] = 16'sd-18;
        fc2_weights[9][21] = 16'sd-45;
        fc2_weights[9][22] = 16'sd-18;
        fc2_weights[9][23] = 16'sd-5;
        fc2_weights[9][24] = 16'sd-51;
        fc2_weights[9][25] = 16'sd59;
        fc2_weights[9][26] = 16'sd-55;
        fc2_weights[9][27] = 16'sd6;
        fc2_weights[9][28] = 16'sd-14;
        fc2_weights[9][29] = 16'sd-10;
        fc2_weights[9][30] = 16'sd-14;
        fc2_weights[9][31] = 16'sd-45;
        fc2_weights[9][32] = 16'sd-50;
        fc2_weights[9][33] = 16'sd-58;
        fc2_weights[9][34] = 16'sd-7;
        fc2_weights[9][35] = 16'sd39;
        fc2_weights[9][36] = 16'sd-13;
        fc2_weights[9][37] = 16'sd-74;
        fc2_weights[9][38] = 16'sd74;
        fc2_weights[9][39] = 16'sd23;
        fc2_weights[9][40] = 16'sd-5;
        fc2_weights[9][41] = 16'sd59;
        fc2_weights[9][42] = 16'sd0;
        fc2_weights[9][43] = 16'sd1;
        fc2_weights[9][44] = 16'sd35;
        fc2_weights[9][45] = 16'sd74;
        fc2_weights[9][46] = 16'sd100;
        fc2_weights[9][47] = 16'sd-40;
        fc2_weights[9][48] = 16'sd22;
        fc2_weights[9][49] = 16'sd13;
        fc2_weights[9][50] = 16'sd13;
        fc2_weights[9][51] = 16'sd-25;
        fc2_weights[9][52] = 16'sd-54;
        fc2_weights[9][53] = 16'sd34;
        fc2_weights[9][54] = 16'sd-27;
        fc2_weights[9][55] = 16'sd34;
        fc2_weights[9][56] = 16'sd54;
        fc2_weights[9][57] = 16'sd12;
        fc2_weights[9][58] = 16'sd26;
        fc2_weights[9][59] = 16'sd-7;
        fc2_weights[9][60] = 16'sd33;
        fc2_weights[9][61] = 16'sd-70;
        fc2_weights[9][62] = 16'sd-20;
        fc2_weights[9][63] = 16'sd38;
        fc2_weights[9][64] = 16'sd-42;
        fc2_weights[9][65] = 16'sd46;
        fc2_weights[9][66] = 16'sd-45;
        fc2_weights[9][67] = 16'sd-10;
        fc2_weights[9][68] = 16'sd-57;
        fc2_weights[9][69] = 16'sd19;
        fc2_weights[9][70] = 16'sd39;
        fc2_weights[9][71] = 16'sd18;
        fc2_weights[9][72] = 16'sd10;
        fc2_weights[9][73] = 16'sd-109;
        fc2_weights[9][74] = 16'sd57;
        fc2_weights[9][75] = 16'sd13;
        fc2_weights[9][76] = 16'sd-58;
        fc2_weights[9][77] = 16'sd51;
        fc2_weights[9][78] = 16'sd-33;
        fc2_weights[9][79] = 16'sd-1;
        fc2_weights[9][80] = 16'sd-77;
        fc2_weights[9][81] = 16'sd0;
        fc2_weights[9][82] = 16'sd0;
        fc2_weights[9][83] = 16'sd-17;
        fc2_weights[9][84] = 16'sd-20;
        fc2_weights[9][85] = 16'sd-23;
        fc2_weights[9][86] = 16'sd-2;
        fc2_weights[9][87] = 16'sd-85;
        fc2_weights[9][88] = 16'sd87;
        fc2_weights[9][89] = 16'sd7;
        fc2_weights[9][90] = 16'sd27;
        fc2_weights[9][91] = 16'sd-13;
        fc2_weights[9][92] = 16'sd47;
        fc2_weights[9][93] = 16'sd-20;
        fc2_weights[9][94] = 16'sd23;
        fc2_weights[9][95] = 16'sd1;
        fc2_weights[9][96] = 16'sd50;
        fc2_weights[9][97] = 16'sd21;
        fc2_weights[9][98] = 16'sd39;
        fc2_weights[9][99] = 16'sd-10;
        fc2_weights[9][100] = 16'sd38;
        fc2_weights[9][101] = 16'sd-13;
        fc2_weights[9][102] = 16'sd49;
        fc2_weights[9][103] = 16'sd13;
        fc2_weights[9][104] = 16'sd107;
        fc2_weights[9][105] = 16'sd-36;
        fc2_weights[9][106] = 16'sd19;
        fc2_weights[9][107] = 16'sd33;
        fc2_weights[9][108] = 16'sd-49;
        fc2_weights[9][109] = 16'sd-49;
        fc2_weights[9][110] = 16'sd60;
        fc2_weights[9][111] = 16'sd23;
        fc2_weights[9][112] = 16'sd-11;
        fc2_weights[9][113] = 16'sd-30;
        fc2_weights[9][114] = 16'sd-29;
        fc2_weights[9][115] = 16'sd-21;
        fc2_weights[9][116] = 16'sd5;
        fc2_weights[9][117] = 16'sd-33;
        fc2_weights[9][118] = 16'sd-2;
        fc2_weights[9][119] = 16'sd-4;
        fc2_weights[9][120] = 16'sd15;
        fc2_weights[9][121] = 16'sd30;
        fc2_weights[9][122] = 16'sd76;
        fc2_weights[9][123] = 16'sd54;
        fc2_weights[9][124] = 16'sd2;
        fc2_weights[9][125] = 16'sd-7;
        fc2_weights[9][126] = 16'sd-11;
        fc2_weights[9][127] = 16'sd-116;
        fc2_weights[10][0] = 16'sd57;
        fc2_weights[10][1] = 16'sd30;
        fc2_weights[10][2] = 16'sd-29;
        fc2_weights[10][3] = 16'sd112;
        fc2_weights[10][4] = 16'sd-17;
        fc2_weights[10][5] = 16'sd1;
        fc2_weights[10][6] = 16'sd26;
        fc2_weights[10][7] = 16'sd-16;
        fc2_weights[10][8] = 16'sd84;
        fc2_weights[10][9] = 16'sd24;
        fc2_weights[10][10] = 16'sd-61;
        fc2_weights[10][11] = 16'sd23;
        fc2_weights[10][12] = 16'sd89;
        fc2_weights[10][13] = 16'sd7;
        fc2_weights[10][14] = 16'sd-62;
        fc2_weights[10][15] = 16'sd-28;
        fc2_weights[10][16] = 16'sd-23;
        fc2_weights[10][17] = 16'sd26;
        fc2_weights[10][18] = 16'sd38;
        fc2_weights[10][19] = 16'sd25;
        fc2_weights[10][20] = 16'sd23;
        fc2_weights[10][21] = 16'sd26;
        fc2_weights[10][22] = 16'sd-22;
        fc2_weights[10][23] = 16'sd-60;
        fc2_weights[10][24] = 16'sd-17;
        fc2_weights[10][25] = 16'sd-21;
        fc2_weights[10][26] = 16'sd-44;
        fc2_weights[10][27] = 16'sd-11;
        fc2_weights[10][28] = 16'sd-2;
        fc2_weights[10][29] = 16'sd-8;
        fc2_weights[10][30] = 16'sd-9;
        fc2_weights[10][31] = 16'sd-3;
        fc2_weights[10][32] = 16'sd-13;
        fc2_weights[10][33] = 16'sd87;
        fc2_weights[10][34] = 16'sd-15;
        fc2_weights[10][35] = 16'sd-54;
        fc2_weights[10][36] = 16'sd16;
        fc2_weights[10][37] = 16'sd-23;
        fc2_weights[10][38] = 16'sd-6;
        fc2_weights[10][39] = 16'sd22;
        fc2_weights[10][40] = 16'sd-1;
        fc2_weights[10][41] = 16'sd-48;
        fc2_weights[10][42] = 16'sd-57;
        fc2_weights[10][43] = 16'sd1;
        fc2_weights[10][44] = 16'sd-5;
        fc2_weights[10][45] = 16'sd-47;
        fc2_weights[10][46] = 16'sd-35;
        fc2_weights[10][47] = 16'sd19;
        fc2_weights[10][48] = 16'sd-55;
        fc2_weights[10][49] = 16'sd-34;
        fc2_weights[10][50] = 16'sd-14;
        fc2_weights[10][51] = 16'sd-62;
        fc2_weights[10][52] = 16'sd-64;
        fc2_weights[10][53] = 16'sd-43;
        fc2_weights[10][54] = 16'sd-11;
        fc2_weights[10][55] = 16'sd-38;
        fc2_weights[10][56] = 16'sd-10;
        fc2_weights[10][57] = 16'sd-38;
        fc2_weights[10][58] = 16'sd-60;
        fc2_weights[10][59] = 16'sd3;
        fc2_weights[10][60] = 16'sd-81;
        fc2_weights[10][61] = 16'sd-10;
        fc2_weights[10][62] = 16'sd-37;
        fc2_weights[10][63] = 16'sd-39;
        fc2_weights[10][64] = 16'sd-23;
        fc2_weights[10][65] = 16'sd-55;
        fc2_weights[10][66] = 16'sd-38;
        fc2_weights[10][67] = 16'sd-9;
        fc2_weights[10][68] = 16'sd68;
        fc2_weights[10][69] = 16'sd4;
        fc2_weights[10][70] = 16'sd-36;
        fc2_weights[10][71] = 16'sd-53;
        fc2_weights[10][72] = 16'sd23;
        fc2_weights[10][73] = 16'sd-8;
        fc2_weights[10][74] = 16'sd-3;
        fc2_weights[10][75] = 16'sd-27;
        fc2_weights[10][76] = 16'sd-23;
        fc2_weights[10][77] = 16'sd17;
        fc2_weights[10][78] = 16'sd63;
        fc2_weights[10][79] = 16'sd20;
        fc2_weights[10][80] = 16'sd68;
        fc2_weights[10][81] = 16'sd-55;
        fc2_weights[10][82] = 16'sd-6;
        fc2_weights[10][83] = 16'sd-37;
        fc2_weights[10][84] = 16'sd43;
        fc2_weights[10][85] = 16'sd-16;
        fc2_weights[10][86] = 16'sd-60;
        fc2_weights[10][87] = 16'sd64;
        fc2_weights[10][88] = 16'sd-29;
        fc2_weights[10][89] = 16'sd-29;
        fc2_weights[10][90] = 16'sd-29;
        fc2_weights[10][91] = 16'sd-11;
        fc2_weights[10][92] = 16'sd-37;
        fc2_weights[10][93] = 16'sd119;
        fc2_weights[10][94] = 16'sd27;
        fc2_weights[10][95] = 16'sd-4;
        fc2_weights[10][96] = 16'sd-85;
        fc2_weights[10][97] = 16'sd-14;
        fc2_weights[10][98] = 16'sd-42;
        fc2_weights[10][99] = 16'sd22;
        fc2_weights[10][100] = 16'sd-110;
        fc2_weights[10][101] = 16'sd52;
        fc2_weights[10][102] = 16'sd-63;
        fc2_weights[10][103] = 16'sd-17;
        fc2_weights[10][104] = 16'sd-11;
        fc2_weights[10][105] = 16'sd-33;
        fc2_weights[10][106] = 16'sd-13;
        fc2_weights[10][107] = 16'sd-68;
        fc2_weights[10][108] = 16'sd-3;
        fc2_weights[10][109] = 16'sd-42;
        fc2_weights[10][110] = 16'sd-4;
        fc2_weights[10][111] = 16'sd-28;
        fc2_weights[10][112] = 16'sd44;
        fc2_weights[10][113] = 16'sd54;
        fc2_weights[10][114] = 16'sd-140;
        fc2_weights[10][115] = 16'sd14;
        fc2_weights[10][116] = 16'sd-2;
        fc2_weights[10][117] = 16'sd28;
        fc2_weights[10][118] = 16'sd32;
        fc2_weights[10][119] = 16'sd-28;
        fc2_weights[10][120] = 16'sd100;
        fc2_weights[10][121] = 16'sd-14;
        fc2_weights[10][122] = 16'sd-81;
        fc2_weights[10][123] = 16'sd-16;
        fc2_weights[10][124] = 16'sd20;
        fc2_weights[10][125] = 16'sd-24;
        fc2_weights[10][126] = 16'sd-34;
        fc2_weights[10][127] = 16'sd-55;
        fc2_weights[11][0] = 16'sd-21;
        fc2_weights[11][1] = 16'sd-7;
        fc2_weights[11][2] = 16'sd-22;
        fc2_weights[11][3] = 16'sd-20;
        fc2_weights[11][4] = 16'sd-46;
        fc2_weights[11][5] = 16'sd-30;
        fc2_weights[11][6] = 16'sd-33;
        fc2_weights[11][7] = 16'sd-30;
        fc2_weights[11][8] = 16'sd-22;
        fc2_weights[11][9] = 16'sd-5;
        fc2_weights[11][10] = 16'sd-5;
        fc2_weights[11][11] = 16'sd-39;
        fc2_weights[11][12] = 16'sd0;
        fc2_weights[11][13] = 16'sd-12;
        fc2_weights[11][14] = 16'sd21;
        fc2_weights[11][15] = 16'sd14;
        fc2_weights[11][16] = 16'sd-39;
        fc2_weights[11][17] = 16'sd-13;
        fc2_weights[11][18] = 16'sd58;
        fc2_weights[11][19] = 16'sd3;
        fc2_weights[11][20] = 16'sd31;
        fc2_weights[11][21] = 16'sd-37;
        fc2_weights[11][22] = 16'sd8;
        fc2_weights[11][23] = 16'sd2;
        fc2_weights[11][24] = 16'sd13;
        fc2_weights[11][25] = 16'sd38;
        fc2_weights[11][26] = 16'sd-20;
        fc2_weights[11][27] = 16'sd6;
        fc2_weights[11][28] = 16'sd-51;
        fc2_weights[11][29] = 16'sd3;
        fc2_weights[11][30] = 16'sd-9;
        fc2_weights[11][31] = 16'sd14;
        fc2_weights[11][32] = 16'sd36;
        fc2_weights[11][33] = 16'sd2;
        fc2_weights[11][34] = 16'sd67;
        fc2_weights[11][35] = 16'sd-17;
        fc2_weights[11][36] = 16'sd-24;
        fc2_weights[11][37] = 16'sd-21;
        fc2_weights[11][38] = 16'sd-11;
        fc2_weights[11][39] = 16'sd-22;
        fc2_weights[11][40] = 16'sd-32;
        fc2_weights[11][41] = 16'sd24;
        fc2_weights[11][42] = 16'sd15;
        fc2_weights[11][43] = 16'sd26;
        fc2_weights[11][44] = 16'sd8;
        fc2_weights[11][45] = 16'sd66;
        fc2_weights[11][46] = 16'sd38;
        fc2_weights[11][47] = 16'sd-8;
        fc2_weights[11][48] = 16'sd26;
        fc2_weights[11][49] = 16'sd-1;
        fc2_weights[11][50] = 16'sd32;
        fc2_weights[11][51] = 16'sd-35;
        fc2_weights[11][52] = 16'sd42;
        fc2_weights[11][53] = 16'sd56;
        fc2_weights[11][54] = 16'sd0;
        fc2_weights[11][55] = 16'sd-12;
        fc2_weights[11][56] = 16'sd-12;
        fc2_weights[11][57] = 16'sd7;
        fc2_weights[11][58] = 16'sd21;
        fc2_weights[11][59] = 16'sd26;
        fc2_weights[11][60] = 16'sd-18;
        fc2_weights[11][61] = 16'sd-53;
        fc2_weights[11][62] = 16'sd9;
        fc2_weights[11][63] = 16'sd42;
        fc2_weights[11][64] = 16'sd-38;
        fc2_weights[11][65] = 16'sd38;
        fc2_weights[11][66] = 16'sd12;
        fc2_weights[11][67] = 16'sd-24;
        fc2_weights[11][68] = 16'sd5;
        fc2_weights[11][69] = 16'sd76;
        fc2_weights[11][70] = 16'sd21;
        fc2_weights[11][71] = 16'sd-37;
        fc2_weights[11][72] = 16'sd15;
        fc2_weights[11][73] = 16'sd-37;
        fc2_weights[11][74] = 16'sd21;
        fc2_weights[11][75] = 16'sd-42;
        fc2_weights[11][76] = 16'sd7;
        fc2_weights[11][77] = 16'sd18;
        fc2_weights[11][78] = 16'sd-44;
        fc2_weights[11][79] = 16'sd-41;
        fc2_weights[11][80] = 16'sd-17;
        fc2_weights[11][81] = 16'sd-29;
        fc2_weights[11][82] = 16'sd-11;
        fc2_weights[11][83] = 16'sd-14;
        fc2_weights[11][84] = 16'sd60;
        fc2_weights[11][85] = 16'sd6;
        fc2_weights[11][86] = 16'sd-32;
        fc2_weights[11][87] = 16'sd-18;
        fc2_weights[11][88] = 16'sd76;
        fc2_weights[11][89] = 16'sd-26;
        fc2_weights[11][90] = 16'sd30;
        fc2_weights[11][91] = 16'sd-18;
        fc2_weights[11][92] = 16'sd26;
        fc2_weights[11][93] = 16'sd-51;
        fc2_weights[11][94] = 16'sd18;
        fc2_weights[11][95] = 16'sd-5;
        fc2_weights[11][96] = 16'sd53;
        fc2_weights[11][97] = 16'sd-20;
        fc2_weights[11][98] = 16'sd-9;
        fc2_weights[11][99] = 16'sd-23;
        fc2_weights[11][100] = 16'sd29;
        fc2_weights[11][101] = 16'sd-19;
        fc2_weights[11][102] = 16'sd30;
        fc2_weights[11][103] = 16'sd9;
        fc2_weights[11][104] = 16'sd5;
        fc2_weights[11][105] = 16'sd-51;
        fc2_weights[11][106] = 16'sd7;
        fc2_weights[11][107] = 16'sd59;
        fc2_weights[11][108] = 16'sd-6;
        fc2_weights[11][109] = 16'sd5;
        fc2_weights[11][110] = 16'sd69;
        fc2_weights[11][111] = 16'sd4;
        fc2_weights[11][112] = 16'sd-30;
        fc2_weights[11][113] = 16'sd-8;
        fc2_weights[11][114] = 16'sd18;
        fc2_weights[11][115] = 16'sd-19;
        fc2_weights[11][116] = 16'sd18;
        fc2_weights[11][117] = 16'sd53;
        fc2_weights[11][118] = 16'sd-2;
        fc2_weights[11][119] = 16'sd-32;
        fc2_weights[11][120] = 16'sd8;
        fc2_weights[11][121] = 16'sd47;
        fc2_weights[11][122] = 16'sd65;
        fc2_weights[11][123] = 16'sd26;
        fc2_weights[11][124] = 16'sd-1;
        fc2_weights[11][125] = 16'sd28;
        fc2_weights[11][126] = 16'sd26;
        fc2_weights[11][127] = 16'sd-6;
        fc2_weights[12][0] = 16'sd-30;
        fc2_weights[12][1] = 16'sd-70;
        fc2_weights[12][2] = 16'sd30;
        fc2_weights[12][3] = 16'sd-48;
        fc2_weights[12][4] = 16'sd-2;
        fc2_weights[12][5] = 16'sd-33;
        fc2_weights[12][6] = 16'sd18;
        fc2_weights[12][7] = 16'sd-1;
        fc2_weights[12][8] = 16'sd16;
        fc2_weights[12][9] = 16'sd-49;
        fc2_weights[12][10] = 16'sd41;
        fc2_weights[12][11] = 16'sd-1;
        fc2_weights[12][12] = 16'sd-22;
        fc2_weights[12][13] = 16'sd-30;
        fc2_weights[12][14] = 16'sd45;
        fc2_weights[12][15] = 16'sd-24;
        fc2_weights[12][16] = 16'sd44;
        fc2_weights[12][17] = 16'sd-88;
        fc2_weights[12][18] = 16'sd-7;
        fc2_weights[12][19] = 16'sd-39;
        fc2_weights[12][20] = 16'sd-78;
        fc2_weights[12][21] = 16'sd55;
        fc2_weights[12][22] = 16'sd26;
        fc2_weights[12][23] = 16'sd60;
        fc2_weights[12][24] = 16'sd-31;
        fc2_weights[12][25] = 16'sd-27;
        fc2_weights[12][26] = 16'sd40;
        fc2_weights[12][27] = 16'sd-2;
        fc2_weights[12][28] = 16'sd-34;
        fc2_weights[12][29] = 16'sd38;
        fc2_weights[12][30] = 16'sd-41;
        fc2_weights[12][31] = 16'sd-12;
        fc2_weights[12][32] = 16'sd-36;
        fc2_weights[12][33] = 16'sd-17;
        fc2_weights[12][34] = 16'sd-61;
        fc2_weights[12][35] = 16'sd27;
        fc2_weights[12][36] = 16'sd12;
        fc2_weights[12][37] = 16'sd-1;
        fc2_weights[12][38] = 16'sd3;
        fc2_weights[12][39] = 16'sd-41;
        fc2_weights[12][40] = 16'sd-22;
        fc2_weights[12][41] = 16'sd17;
        fc2_weights[12][42] = 16'sd-11;
        fc2_weights[12][43] = 16'sd-60;
        fc2_weights[12][44] = 16'sd-47;
        fc2_weights[12][45] = 16'sd89;
        fc2_weights[12][46] = 16'sd29;
        fc2_weights[12][47] = 16'sd13;
        fc2_weights[12][48] = 16'sd-13;
        fc2_weights[12][49] = 16'sd13;
        fc2_weights[12][50] = 16'sd-52;
        fc2_weights[12][51] = 16'sd63;
        fc2_weights[12][52] = 16'sd-44;
        fc2_weights[12][53] = 16'sd16;
        fc2_weights[12][54] = 16'sd121;
        fc2_weights[12][55] = 16'sd27;
        fc2_weights[12][56] = 16'sd-7;
        fc2_weights[12][57] = 16'sd-9;
        fc2_weights[12][58] = 16'sd-17;
        fc2_weights[12][59] = 16'sd-60;
        fc2_weights[12][60] = 16'sd47;
        fc2_weights[12][61] = 16'sd36;
        fc2_weights[12][62] = 16'sd32;
        fc2_weights[12][63] = 16'sd4;
        fc2_weights[12][64] = 16'sd25;
        fc2_weights[12][65] = 16'sd-4;
        fc2_weights[12][66] = 16'sd36;
        fc2_weights[12][67] = 16'sd17;
        fc2_weights[12][68] = 16'sd-50;
        fc2_weights[12][69] = 16'sd2;
        fc2_weights[12][70] = 16'sd17;
        fc2_weights[12][71] = 16'sd6;
        fc2_weights[12][72] = 16'sd-28;
        fc2_weights[12][73] = 16'sd-63;
        fc2_weights[12][74] = 16'sd-19;
        fc2_weights[12][75] = 16'sd14;
        fc2_weights[12][76] = 16'sd9;
        fc2_weights[12][77] = 16'sd33;
        fc2_weights[12][78] = 16'sd-37;
        fc2_weights[12][79] = 16'sd-7;
        fc2_weights[12][80] = 16'sd4;
        fc2_weights[12][81] = 16'sd24;
        fc2_weights[12][82] = 16'sd13;
        fc2_weights[12][83] = 16'sd23;
        fc2_weights[12][84] = 16'sd-27;
        fc2_weights[12][85] = 16'sd10;
        fc2_weights[12][86] = 16'sd-6;
        fc2_weights[12][87] = 16'sd-58;
        fc2_weights[12][88] = 16'sd3;
        fc2_weights[12][89] = 16'sd9;
        fc2_weights[12][90] = 16'sd-9;
        fc2_weights[12][91] = 16'sd74;
        fc2_weights[12][92] = 16'sd-16;
        fc2_weights[12][93] = 16'sd-18;
        fc2_weights[12][94] = 16'sd-42;
        fc2_weights[12][95] = 16'sd54;
        fc2_weights[12][96] = 16'sd-63;
        fc2_weights[12][97] = 16'sd-16;
        fc2_weights[12][98] = 16'sd76;
        fc2_weights[12][99] = 16'sd-21;
        fc2_weights[12][100] = 16'sd33;
        fc2_weights[12][101] = 16'sd-26;
        fc2_weights[12][102] = 16'sd50;
        fc2_weights[12][103] = 16'sd36;
        fc2_weights[12][104] = 16'sd41;
        fc2_weights[12][105] = 16'sd-33;
        fc2_weights[12][106] = 16'sd4;
        fc2_weights[12][107] = 16'sd-17;
        fc2_weights[12][108] = 16'sd-11;
        fc2_weights[12][109] = 16'sd-13;
        fc2_weights[12][110] = 16'sd-18;
        fc2_weights[12][111] = 16'sd19;
        fc2_weights[12][112] = 16'sd-15;
        fc2_weights[12][113] = 16'sd-25;
        fc2_weights[12][114] = 16'sd10;
        fc2_weights[12][115] = 16'sd-2;
        fc2_weights[12][116] = 16'sd37;
        fc2_weights[12][117] = 16'sd-46;
        fc2_weights[12][118] = 16'sd15;
        fc2_weights[12][119] = 16'sd-36;
        fc2_weights[12][120] = 16'sd-44;
        fc2_weights[12][121] = 16'sd15;
        fc2_weights[12][122] = 16'sd-9;
        fc2_weights[12][123] = 16'sd13;
        fc2_weights[12][124] = 16'sd-45;
        fc2_weights[12][125] = 16'sd9;
        fc2_weights[12][126] = 16'sd3;
        fc2_weights[12][127] = 16'sd10;
        fc2_weights[13][0] = 16'sd-7;
        fc2_weights[13][1] = 16'sd-46;
        fc2_weights[13][2] = 16'sd25;
        fc2_weights[13][3] = 16'sd-11;
        fc2_weights[13][4] = 16'sd-3;
        fc2_weights[13][5] = 16'sd-34;
        fc2_weights[13][6] = 16'sd-15;
        fc2_weights[13][7] = 16'sd36;
        fc2_weights[13][8] = 16'sd-44;
        fc2_weights[13][9] = 16'sd56;
        fc2_weights[13][10] = 16'sd14;
        fc2_weights[13][11] = 16'sd-18;
        fc2_weights[13][12] = 16'sd5;
        fc2_weights[13][13] = 16'sd-16;
        fc2_weights[13][14] = 16'sd-18;
        fc2_weights[13][15] = 16'sd16;
        fc2_weights[13][16] = 16'sd-12;
        fc2_weights[13][17] = 16'sd-33;
        fc2_weights[13][18] = 16'sd11;
        fc2_weights[13][19] = 16'sd-13;
        fc2_weights[13][20] = 16'sd-24;
        fc2_weights[13][21] = 16'sd-33;
        fc2_weights[13][22] = 16'sd79;
        fc2_weights[13][23] = 16'sd-21;
        fc2_weights[13][24] = 16'sd-20;
        fc2_weights[13][25] = 16'sd-16;
        fc2_weights[13][26] = 16'sd0;
        fc2_weights[13][27] = 16'sd7;
        fc2_weights[13][28] = 16'sd-10;
        fc2_weights[13][29] = 16'sd39;
        fc2_weights[13][30] = 16'sd2;
        fc2_weights[13][31] = 16'sd0;
        fc2_weights[13][32] = 16'sd3;
        fc2_weights[13][33] = 16'sd57;
        fc2_weights[13][34] = 16'sd16;
        fc2_weights[13][35] = 16'sd9;
        fc2_weights[13][36] = 16'sd1;
        fc2_weights[13][37] = 16'sd27;
        fc2_weights[13][38] = 16'sd25;
        fc2_weights[13][39] = 16'sd49;
        fc2_weights[13][40] = 16'sd-25;
        fc2_weights[13][41] = 16'sd-9;
        fc2_weights[13][42] = 16'sd27;
        fc2_weights[13][43] = 16'sd77;
        fc2_weights[13][44] = 16'sd-30;
        fc2_weights[13][45] = 16'sd-42;
        fc2_weights[13][46] = 16'sd-22;
        fc2_weights[13][47] = 16'sd-9;
        fc2_weights[13][48] = 16'sd-12;
        fc2_weights[13][49] = 16'sd-18;
        fc2_weights[13][50] = 16'sd16;
        fc2_weights[13][51] = 16'sd21;
        fc2_weights[13][52] = 16'sd46;
        fc2_weights[13][53] = 16'sd30;
        fc2_weights[13][54] = 16'sd30;
        fc2_weights[13][55] = 16'sd-32;
        fc2_weights[13][56] = 16'sd16;
        fc2_weights[13][57] = 16'sd-34;
        fc2_weights[13][58] = 16'sd6;
        fc2_weights[13][59] = 16'sd-36;
        fc2_weights[13][60] = 16'sd-35;
        fc2_weights[13][61] = 16'sd1;
        fc2_weights[13][62] = 16'sd44;
        fc2_weights[13][63] = 16'sd-21;
        fc2_weights[13][64] = 16'sd-20;
        fc2_weights[13][65] = 16'sd-9;
        fc2_weights[13][66] = 16'sd-37;
        fc2_weights[13][67] = 16'sd-1;
        fc2_weights[13][68] = 16'sd28;
        fc2_weights[13][69] = 16'sd-52;
        fc2_weights[13][70] = 16'sd-22;
        fc2_weights[13][71] = 16'sd23;
        fc2_weights[13][72] = 16'sd-21;
        fc2_weights[13][73] = 16'sd-24;
        fc2_weights[13][74] = 16'sd45;
        fc2_weights[13][75] = 16'sd28;
        fc2_weights[13][76] = 16'sd-20;
        fc2_weights[13][77] = 16'sd17;
        fc2_weights[13][78] = 16'sd-30;
        fc2_weights[13][79] = 16'sd-30;
        fc2_weights[13][80] = 16'sd-26;
        fc2_weights[13][81] = 16'sd8;
        fc2_weights[13][82] = 16'sd50;
        fc2_weights[13][83] = 16'sd3;
        fc2_weights[13][84] = 16'sd-12;
        fc2_weights[13][85] = 16'sd-3;
        fc2_weights[13][86] = 16'sd-10;
        fc2_weights[13][87] = 16'sd-32;
        fc2_weights[13][88] = 16'sd-35;
        fc2_weights[13][89] = 16'sd-25;
        fc2_weights[13][90] = 16'sd28;
        fc2_weights[13][91] = 16'sd-28;
        fc2_weights[13][92] = 16'sd-21;
        fc2_weights[13][93] = 16'sd25;
        fc2_weights[13][94] = 16'sd53;
        fc2_weights[13][95] = 16'sd21;
        fc2_weights[13][96] = 16'sd-19;
        fc2_weights[13][97] = 16'sd57;
        fc2_weights[13][98] = 16'sd17;
        fc2_weights[13][99] = 16'sd12;
        fc2_weights[13][100] = 16'sd-29;
        fc2_weights[13][101] = 16'sd3;
        fc2_weights[13][102] = 16'sd-30;
        fc2_weights[13][103] = 16'sd17;
        fc2_weights[13][104] = 16'sd-31;
        fc2_weights[13][105] = 16'sd3;
        fc2_weights[13][106] = 16'sd22;
        fc2_weights[13][107] = 16'sd-25;
        fc2_weights[13][108] = 16'sd18;
        fc2_weights[13][109] = 16'sd-10;
        fc2_weights[13][110] = 16'sd-14;
        fc2_weights[13][111] = 16'sd20;
        fc2_weights[13][112] = 16'sd41;
        fc2_weights[13][113] = 16'sd5;
        fc2_weights[13][114] = 16'sd-16;
        fc2_weights[13][115] = 16'sd-25;
        fc2_weights[13][116] = 16'sd19;
        fc2_weights[13][117] = 16'sd-28;
        fc2_weights[13][118] = 16'sd6;
        fc2_weights[13][119] = 16'sd-29;
        fc2_weights[13][120] = 16'sd-25;
        fc2_weights[13][121] = 16'sd8;
        fc2_weights[13][122] = 16'sd6;
        fc2_weights[13][123] = 16'sd-8;
        fc2_weights[13][124] = 16'sd18;
        fc2_weights[13][125] = 16'sd11;
        fc2_weights[13][126] = 16'sd-10;
        fc2_weights[13][127] = 16'sd-18;
        fc2_weights[14][0] = 16'sd-4;
        fc2_weights[14][1] = 16'sd-25;
        fc2_weights[14][2] = 16'sd96;
        fc2_weights[14][3] = 16'sd-71;
        fc2_weights[14][4] = 16'sd-13;
        fc2_weights[14][5] = 16'sd-34;
        fc2_weights[14][6] = 16'sd-42;
        fc2_weights[14][7] = 16'sd15;
        fc2_weights[14][8] = 16'sd-27;
        fc2_weights[14][9] = 16'sd-56;
        fc2_weights[14][10] = 16'sd8;
        fc2_weights[14][11] = 16'sd-41;
        fc2_weights[14][12] = 16'sd-4;
        fc2_weights[14][13] = 16'sd-30;
        fc2_weights[14][14] = 16'sd13;
        fc2_weights[14][15] = 16'sd31;
        fc2_weights[14][16] = 16'sd-2;
        fc2_weights[14][17] = 16'sd-42;
        fc2_weights[14][18] = 16'sd18;
        fc2_weights[14][19] = 16'sd-28;
        fc2_weights[14][20] = 16'sd34;
        fc2_weights[14][21] = 16'sd-55;
        fc2_weights[14][22] = 16'sd-9;
        fc2_weights[14][23] = 16'sd10;
        fc2_weights[14][24] = 16'sd-4;
        fc2_weights[14][25] = 16'sd25;
        fc2_weights[14][26] = 16'sd19;
        fc2_weights[14][27] = 16'sd-3;
        fc2_weights[14][28] = 16'sd-80;
        fc2_weights[14][29] = 16'sd-21;
        fc2_weights[14][30] = 16'sd-27;
        fc2_weights[14][31] = 16'sd24;
        fc2_weights[14][32] = 16'sd-14;
        fc2_weights[14][33] = 16'sd-38;
        fc2_weights[14][34] = 16'sd53;
        fc2_weights[14][35] = 16'sd17;
        fc2_weights[14][36] = 16'sd41;
        fc2_weights[14][37] = 16'sd-87;
        fc2_weights[14][38] = 16'sd44;
        fc2_weights[14][39] = 16'sd-54;
        fc2_weights[14][40] = 16'sd-93;
        fc2_weights[14][41] = 16'sd72;
        fc2_weights[14][42] = 16'sd-45;
        fc2_weights[14][43] = 16'sd-1;
        fc2_weights[14][44] = 16'sd20;
        fc2_weights[14][45] = 16'sd94;
        fc2_weights[14][46] = 16'sd23;
        fc2_weights[14][47] = 16'sd-16;
        fc2_weights[14][48] = 16'sd13;
        fc2_weights[14][49] = 16'sd70;
        fc2_weights[14][50] = 16'sd9;
        fc2_weights[14][51] = 16'sd-39;
        fc2_weights[14][52] = 16'sd24;
        fc2_weights[14][53] = 16'sd-36;
        fc2_weights[14][54] = 16'sd61;
        fc2_weights[14][55] = 16'sd19;
        fc2_weights[14][56] = 16'sd-44;
        fc2_weights[14][57] = 16'sd12;
        fc2_weights[14][58] = 16'sd29;
        fc2_weights[14][59] = 16'sd29;
        fc2_weights[14][60] = 16'sd2;
        fc2_weights[14][61] = 16'sd-39;
        fc2_weights[14][62] = 16'sd-10;
        fc2_weights[14][63] = 16'sd87;
        fc2_weights[14][64] = 16'sd12;
        fc2_weights[14][65] = 16'sd8;
        fc2_weights[14][66] = 16'sd74;
        fc2_weights[14][67] = 16'sd-40;
        fc2_weights[14][68] = 16'sd-23;
        fc2_weights[14][69] = 16'sd-10;
        fc2_weights[14][70] = 16'sd33;
        fc2_weights[14][71] = 16'sd30;
        fc2_weights[14][72] = 16'sd-36;
        fc2_weights[14][73] = 16'sd-98;
        fc2_weights[14][74] = 16'sd2;
        fc2_weights[14][75] = 16'sd-26;
        fc2_weights[14][76] = 16'sd-49;
        fc2_weights[14][77] = 16'sd50;
        fc2_weights[14][78] = 16'sd-18;
        fc2_weights[14][79] = 16'sd-17;
        fc2_weights[14][80] = 16'sd-9;
        fc2_weights[14][81] = 16'sd-7;
        fc2_weights[14][82] = 16'sd-12;
        fc2_weights[14][83] = 16'sd7;
        fc2_weights[14][84] = 16'sd10;
        fc2_weights[14][85] = 16'sd10;
        fc2_weights[14][86] = 16'sd-25;
        fc2_weights[14][87] = 16'sd-25;
        fc2_weights[14][88] = 16'sd26;
        fc2_weights[14][89] = 16'sd-18;
        fc2_weights[14][90] = 16'sd47;
        fc2_weights[14][91] = 16'sd-21;
        fc2_weights[14][92] = 16'sd70;
        fc2_weights[14][93] = 16'sd-17;
        fc2_weights[14][94] = 16'sd-17;
        fc2_weights[14][95] = 16'sd9;
        fc2_weights[14][96] = 16'sd7;
        fc2_weights[14][97] = 16'sd25;
        fc2_weights[14][98] = 16'sd-5;
        fc2_weights[14][99] = 16'sd-6;
        fc2_weights[14][100] = 16'sd65;
        fc2_weights[14][101] = 16'sd-23;
        fc2_weights[14][102] = 16'sd38;
        fc2_weights[14][103] = 16'sd-40;
        fc2_weights[14][104] = 16'sd17;
        fc2_weights[14][105] = 16'sd-31;
        fc2_weights[14][106] = 16'sd-18;
        fc2_weights[14][107] = 16'sd34;
        fc2_weights[14][108] = 16'sd-60;
        fc2_weights[14][109] = 16'sd31;
        fc2_weights[14][110] = 16'sd7;
        fc2_weights[14][111] = 16'sd33;
        fc2_weights[14][112] = 16'sd-50;
        fc2_weights[14][113] = 16'sd-78;
        fc2_weights[14][114] = 16'sd19;
        fc2_weights[14][115] = 16'sd-37;
        fc2_weights[14][116] = 16'sd-8;
        fc2_weights[14][117] = 16'sd-17;
        fc2_weights[14][118] = 16'sd-25;
        fc2_weights[14][119] = 16'sd-33;
        fc2_weights[14][120] = 16'sd-26;
        fc2_weights[14][121] = 16'sd33;
        fc2_weights[14][122] = 16'sd-10;
        fc2_weights[14][123] = 16'sd12;
        fc2_weights[14][124] = 16'sd-4;
        fc2_weights[14][125] = 16'sd25;
        fc2_weights[14][126] = 16'sd2;
        fc2_weights[14][127] = 16'sd-13;
        fc2_weights[15][0] = 16'sd130;
        fc2_weights[15][1] = 16'sd-21;
        fc2_weights[15][2] = 16'sd-62;
        fc2_weights[15][3] = 16'sd4;
        fc2_weights[15][4] = 16'sd-23;
        fc2_weights[15][5] = 16'sd28;
        fc2_weights[15][6] = 16'sd-2;
        fc2_weights[15][7] = 16'sd-36;
        fc2_weights[15][8] = 16'sd-36;
        fc2_weights[15][9] = 16'sd-29;
        fc2_weights[15][10] = 16'sd-22;
        fc2_weights[15][11] = 16'sd13;
        fc2_weights[15][12] = 16'sd-23;
        fc2_weights[15][13] = 16'sd23;
        fc2_weights[15][14] = 16'sd-39;
        fc2_weights[15][15] = 16'sd3;
        fc2_weights[15][16] = 16'sd72;
        fc2_weights[15][17] = 16'sd-22;
        fc2_weights[15][18] = 16'sd1;
        fc2_weights[15][19] = 16'sd12;
        fc2_weights[15][20] = 16'sd-58;
        fc2_weights[15][21] = 16'sd-30;
        fc2_weights[15][22] = 16'sd-54;
        fc2_weights[15][23] = 16'sd-9;
        fc2_weights[15][24] = 16'sd-87;
        fc2_weights[15][25] = 16'sd-8;
        fc2_weights[15][26] = 16'sd-20;
        fc2_weights[15][27] = 16'sd-72;
        fc2_weights[15][28] = 16'sd40;
        fc2_weights[15][29] = 16'sd-37;
        fc2_weights[15][30] = 16'sd18;
        fc2_weights[15][31] = 16'sd20;
        fc2_weights[15][32] = 16'sd-82;
        fc2_weights[15][33] = 16'sd-66;
        fc2_weights[15][34] = 16'sd-36;
        fc2_weights[15][35] = 16'sd49;
        fc2_weights[15][36] = 16'sd-24;
        fc2_weights[15][37] = 16'sd-49;
        fc2_weights[15][38] = 16'sd27;
        fc2_weights[15][39] = 16'sd40;
        fc2_weights[15][40] = 16'sd18;
        fc2_weights[15][41] = 16'sd41;
        fc2_weights[15][42] = 16'sd-47;
        fc2_weights[15][43] = 16'sd-33;
        fc2_weights[15][44] = 16'sd-46;
        fc2_weights[15][45] = 16'sd-21;
        fc2_weights[15][46] = 16'sd-5;
        fc2_weights[15][47] = 16'sd-28;
        fc2_weights[15][48] = 16'sd-56;
        fc2_weights[15][49] = 16'sd4;
        fc2_weights[15][50] = 16'sd-33;
        fc2_weights[15][51] = 16'sd14;
        fc2_weights[15][52] = 16'sd-52;
        fc2_weights[15][53] = 16'sd6;
        fc2_weights[15][54] = 16'sd-34;
        fc2_weights[15][55] = 16'sd19;
        fc2_weights[15][56] = 16'sd56;
        fc2_weights[15][57] = 16'sd-63;
        fc2_weights[15][58] = 16'sd-57;
        fc2_weights[15][59] = 16'sd-45;
        fc2_weights[15][60] = 16'sd-1;
        fc2_weights[15][61] = 16'sd49;
        fc2_weights[15][62] = 16'sd-6;
        fc2_weights[15][63] = 16'sd-27;
        fc2_weights[15][64] = 16'sd10;
        fc2_weights[15][65] = 16'sd20;
        fc2_weights[15][66] = 16'sd-18;
        fc2_weights[15][67] = 16'sd-28;
        fc2_weights[15][68] = 16'sd-25;
        fc2_weights[15][69] = 16'sd13;
        fc2_weights[15][70] = 16'sd48;
        fc2_weights[15][71] = 16'sd3;
        fc2_weights[15][72] = 16'sd61;
        fc2_weights[15][73] = 16'sd-3;
        fc2_weights[15][74] = 16'sd-22;
        fc2_weights[15][75] = 16'sd-12;
        fc2_weights[15][76] = 16'sd-10;
        fc2_weights[15][77] = 16'sd-8;
        fc2_weights[15][78] = 16'sd8;
        fc2_weights[15][79] = 16'sd-43;
        fc2_weights[15][80] = 16'sd26;
        fc2_weights[15][81] = 16'sd-62;
        fc2_weights[15][82] = 16'sd11;
        fc2_weights[15][83] = 16'sd101;
        fc2_weights[15][84] = 16'sd-67;
        fc2_weights[15][85] = 16'sd17;
        fc2_weights[15][86] = 16'sd8;
        fc2_weights[15][87] = 16'sd-73;
        fc2_weights[15][88] = 16'sd-59;
        fc2_weights[15][89] = 16'sd45;
        fc2_weights[15][90] = 16'sd-20;
        fc2_weights[15][91] = 16'sd54;
        fc2_weights[15][92] = 16'sd-39;
        fc2_weights[15][93] = 16'sd-12;
        fc2_weights[15][94] = 16'sd-81;
        fc2_weights[15][95] = 16'sd-38;
        fc2_weights[15][96] = 16'sd65;
        fc2_weights[15][97] = 16'sd-17;
        fc2_weights[15][98] = 16'sd92;
        fc2_weights[15][99] = 16'sd-7;
        fc2_weights[15][100] = 16'sd-41;
        fc2_weights[15][101] = 16'sd60;
        fc2_weights[15][102] = 16'sd-7;
        fc2_weights[15][103] = 16'sd-56;
        fc2_weights[15][104] = 16'sd3;
        fc2_weights[15][105] = 16'sd31;
        fc2_weights[15][106] = 16'sd38;
        fc2_weights[15][107] = 16'sd12;
        fc2_weights[15][108] = 16'sd-50;
        fc2_weights[15][109] = 16'sd-7;
        fc2_weights[15][110] = 16'sd-3;
        fc2_weights[15][111] = 16'sd-33;
        fc2_weights[15][112] = 16'sd17;
        fc2_weights[15][113] = 16'sd48;
        fc2_weights[15][114] = 16'sd27;
        fc2_weights[15][115] = 16'sd37;
        fc2_weights[15][116] = 16'sd11;
        fc2_weights[15][117] = 16'sd-18;
        fc2_weights[15][118] = 16'sd-1;
        fc2_weights[15][119] = 16'sd33;
        fc2_weights[15][120] = 16'sd-9;
        fc2_weights[15][121] = 16'sd0;
        fc2_weights[15][122] = 16'sd-52;
        fc2_weights[15][123] = 16'sd25;
        fc2_weights[15][124] = 16'sd0;
        fc2_weights[15][125] = 16'sd-61;
        fc2_weights[15][126] = 16'sd-5;
        fc2_weights[15][127] = 16'sd-49;
        fc2_weights[16][0] = 16'sd-17;
        fc2_weights[16][1] = 16'sd-26;
        fc2_weights[16][2] = 16'sd17;
        fc2_weights[16][3] = 16'sd-39;
        fc2_weights[16][4] = 16'sd-3;
        fc2_weights[16][5] = 16'sd11;
        fc2_weights[16][6] = 16'sd13;
        fc2_weights[16][7] = 16'sd-13;
        fc2_weights[16][8] = 16'sd-4;
        fc2_weights[16][9] = 16'sd-43;
        fc2_weights[16][10] = 16'sd12;
        fc2_weights[16][11] = 16'sd-27;
        fc2_weights[16][12] = 16'sd-27;
        fc2_weights[16][13] = 16'sd-8;
        fc2_weights[16][14] = 16'sd42;
        fc2_weights[16][15] = 16'sd37;
        fc2_weights[16][16] = 16'sd45;
        fc2_weights[16][17] = 16'sd-51;
        fc2_weights[16][18] = 16'sd10;
        fc2_weights[16][19] = 16'sd-35;
        fc2_weights[16][20] = 16'sd6;
        fc2_weights[16][21] = 16'sd4;
        fc2_weights[16][22] = 16'sd8;
        fc2_weights[16][23] = 16'sd-34;
        fc2_weights[16][24] = 16'sd34;
        fc2_weights[16][25] = 16'sd-35;
        fc2_weights[16][26] = 16'sd16;
        fc2_weights[16][27] = 16'sd-2;
        fc2_weights[16][28] = 16'sd-1;
        fc2_weights[16][29] = 16'sd-28;
        fc2_weights[16][30] = 16'sd-30;
        fc2_weights[16][31] = 16'sd-9;
        fc2_weights[16][32] = 16'sd9;
        fc2_weights[16][33] = 16'sd-27;
        fc2_weights[16][34] = 16'sd-5;
        fc2_weights[16][35] = 16'sd-35;
        fc2_weights[16][36] = 16'sd-15;
        fc2_weights[16][37] = 16'sd-21;
        fc2_weights[16][38] = 16'sd51;
        fc2_weights[16][39] = 16'sd31;
        fc2_weights[16][40] = 16'sd-9;
        fc2_weights[16][41] = 16'sd72;
        fc2_weights[16][42] = 16'sd-12;
        fc2_weights[16][43] = 16'sd-27;
        fc2_weights[16][44] = 16'sd-25;
        fc2_weights[16][45] = 16'sd7;
        fc2_weights[16][46] = 16'sd81;
        fc2_weights[16][47] = 16'sd24;
        fc2_weights[16][48] = 16'sd26;
        fc2_weights[16][49] = 16'sd15;
        fc2_weights[16][50] = 16'sd14;
        fc2_weights[16][51] = 16'sd55;
        fc2_weights[16][52] = 16'sd-4;
        fc2_weights[16][53] = 16'sd-8;
        fc2_weights[16][54] = 16'sd96;
        fc2_weights[16][55] = 16'sd13;
        fc2_weights[16][56] = 16'sd5;
        fc2_weights[16][57] = 16'sd56;
        fc2_weights[16][58] = 16'sd-9;
        fc2_weights[16][59] = 16'sd2;
        fc2_weights[16][60] = 16'sd24;
        fc2_weights[16][61] = 16'sd-24;
        fc2_weights[16][62] = 16'sd-39;
        fc2_weights[16][63] = 16'sd63;
        fc2_weights[16][64] = 16'sd-4;
        fc2_weights[16][65] = 16'sd27;
        fc2_weights[16][66] = 16'sd64;
        fc2_weights[16][67] = 16'sd-38;
        fc2_weights[16][68] = 16'sd4;
        fc2_weights[16][69] = 16'sd-43;
        fc2_weights[16][70] = 16'sd7;
        fc2_weights[16][71] = 16'sd-7;
        fc2_weights[16][72] = 16'sd-42;
        fc2_weights[16][73] = 16'sd-1;
        fc2_weights[16][74] = 16'sd2;
        fc2_weights[16][75] = 16'sd-3;
        fc2_weights[16][76] = 16'sd35;
        fc2_weights[16][77] = 16'sd83;
        fc2_weights[16][78] = 16'sd-51;
        fc2_weights[16][79] = 16'sd31;
        fc2_weights[16][80] = 16'sd3;
        fc2_weights[16][81] = 16'sd27;
        fc2_weights[16][82] = 16'sd-20;
        fc2_weights[16][83] = 16'sd2;
        fc2_weights[16][84] = 16'sd31;
        fc2_weights[16][85] = 16'sd21;
        fc2_weights[16][86] = 16'sd33;
        fc2_weights[16][87] = 16'sd4;
        fc2_weights[16][88] = 16'sd1;
        fc2_weights[16][89] = 16'sd-6;
        fc2_weights[16][90] = 16'sd21;
        fc2_weights[16][91] = 16'sd-36;
        fc2_weights[16][92] = 16'sd33;
        fc2_weights[16][93] = 16'sd30;
        fc2_weights[16][94] = 16'sd-78;
        fc2_weights[16][95] = 16'sd17;
        fc2_weights[16][96] = 16'sd-20;
        fc2_weights[16][97] = 16'sd38;
        fc2_weights[16][98] = 16'sd1;
        fc2_weights[16][99] = 16'sd-11;
        fc2_weights[16][100] = 16'sd31;
        fc2_weights[16][101] = 16'sd6;
        fc2_weights[16][102] = 16'sd-31;
        fc2_weights[16][103] = 16'sd-4;
        fc2_weights[16][104] = 16'sd-33;
        fc2_weights[16][105] = 16'sd-7;
        fc2_weights[16][106] = 16'sd5;
        fc2_weights[16][107] = 16'sd66;
        fc2_weights[16][108] = 16'sd-49;
        fc2_weights[16][109] = 16'sd32;
        fc2_weights[16][110] = 16'sd-22;
        fc2_weights[16][111] = 16'sd13;
        fc2_weights[16][112] = 16'sd-17;
        fc2_weights[16][113] = 16'sd8;
        fc2_weights[16][114] = 16'sd-5;
        fc2_weights[16][115] = 16'sd-5;
        fc2_weights[16][116] = 16'sd31;
        fc2_weights[16][117] = 16'sd3;
        fc2_weights[16][118] = 16'sd-12;
        fc2_weights[16][119] = 16'sd12;
        fc2_weights[16][120] = 16'sd-42;
        fc2_weights[16][121] = 16'sd50;
        fc2_weights[16][122] = 16'sd51;
        fc2_weights[16][123] = 16'sd-9;
        fc2_weights[16][124] = 16'sd22;
        fc2_weights[16][125] = 16'sd-6;
        fc2_weights[16][126] = 16'sd30;
        fc2_weights[16][127] = 16'sd29;
        fc2_weights[17][0] = 16'sd21;
        fc2_weights[17][1] = 16'sd-18;
        fc2_weights[17][2] = 16'sd38;
        fc2_weights[17][3] = 16'sd39;
        fc2_weights[17][4] = 16'sd-45;
        fc2_weights[17][5] = 16'sd-6;
        fc2_weights[17][6] = 16'sd-74;
        fc2_weights[17][7] = 16'sd30;
        fc2_weights[17][8] = 16'sd-60;
        fc2_weights[17][9] = 16'sd2;
        fc2_weights[17][10] = 16'sd-11;
        fc2_weights[17][11] = 16'sd-35;
        fc2_weights[17][12] = 16'sd-28;
        fc2_weights[17][13] = 16'sd28;
        fc2_weights[17][14] = 16'sd14;
        fc2_weights[17][15] = 16'sd25;
        fc2_weights[17][16] = 16'sd-22;
        fc2_weights[17][17] = 16'sd-7;
        fc2_weights[17][18] = 16'sd-5;
        fc2_weights[17][19] = 16'sd-4;
        fc2_weights[17][20] = 16'sd10;
        fc2_weights[17][21] = 16'sd7;
        fc2_weights[17][22] = 16'sd-26;
        fc2_weights[17][23] = 16'sd-14;
        fc2_weights[17][24] = 16'sd-8;
        fc2_weights[17][25] = 16'sd14;
        fc2_weights[17][26] = 16'sd8;
        fc2_weights[17][27] = 16'sd14;
        fc2_weights[17][28] = 16'sd-21;
        fc2_weights[17][29] = 16'sd-39;
        fc2_weights[17][30] = 16'sd-13;
        fc2_weights[17][31] = 16'sd-3;
        fc2_weights[17][32] = 16'sd-12;
        fc2_weights[17][33] = 16'sd-13;
        fc2_weights[17][34] = 16'sd26;
        fc2_weights[17][35] = 16'sd27;
        fc2_weights[17][36] = 16'sd3;
        fc2_weights[17][37] = 16'sd-6;
        fc2_weights[17][38] = 16'sd-8;
        fc2_weights[17][39] = 16'sd-57;
        fc2_weights[17][40] = 16'sd8;
        fc2_weights[17][41] = 16'sd-57;
        fc2_weights[17][42] = 16'sd15;
        fc2_weights[17][43] = 16'sd-11;
        fc2_weights[17][44] = 16'sd68;
        fc2_weights[17][45] = 16'sd75;
        fc2_weights[17][46] = 16'sd41;
        fc2_weights[17][47] = 16'sd-43;
        fc2_weights[17][48] = 16'sd-12;
        fc2_weights[17][49] = 16'sd18;
        fc2_weights[17][50] = 16'sd-23;
        fc2_weights[17][51] = 16'sd-32;
        fc2_weights[17][52] = 16'sd30;
        fc2_weights[17][53] = 16'sd-14;
        fc2_weights[17][54] = 16'sd5;
        fc2_weights[17][55] = 16'sd-49;
        fc2_weights[17][56] = 16'sd-1;
        fc2_weights[17][57] = 16'sd34;
        fc2_weights[17][58] = 16'sd38;
        fc2_weights[17][59] = 16'sd24;
        fc2_weights[17][60] = 16'sd-39;
        fc2_weights[17][61] = 16'sd-60;
        fc2_weights[17][62] = 16'sd20;
        fc2_weights[17][63] = 16'sd55;
        fc2_weights[17][64] = 16'sd-3;
        fc2_weights[17][65] = 16'sd49;
        fc2_weights[17][66] = 16'sd35;
        fc2_weights[17][67] = 16'sd9;
        fc2_weights[17][68] = 16'sd23;
        fc2_weights[17][69] = 16'sd67;
        fc2_weights[17][70] = 16'sd3;
        fc2_weights[17][71] = 16'sd-7;
        fc2_weights[17][72] = 16'sd-22;
        fc2_weights[17][73] = 16'sd-24;
        fc2_weights[17][74] = 16'sd42;
        fc2_weights[17][75] = 16'sd-38;
        fc2_weights[17][76] = 16'sd-12;
        fc2_weights[17][77] = 16'sd-23;
        fc2_weights[17][78] = 16'sd-11;
        fc2_weights[17][79] = 16'sd-5;
        fc2_weights[17][80] = 16'sd-71;
        fc2_weights[17][81] = 16'sd17;
        fc2_weights[17][82] = 16'sd-18;
        fc2_weights[17][83] = 16'sd25;
        fc2_weights[17][84] = 16'sd10;
        fc2_weights[17][85] = 16'sd-57;
        fc2_weights[17][86] = 16'sd-1;
        fc2_weights[17][87] = 16'sd-2;
        fc2_weights[17][88] = 16'sd9;
        fc2_weights[17][89] = 16'sd-16;
        fc2_weights[17][90] = 16'sd66;
        fc2_weights[17][91] = 16'sd-34;
        fc2_weights[17][92] = 16'sd12;
        fc2_weights[17][93] = 16'sd-51;
        fc2_weights[17][94] = 16'sd92;
        fc2_weights[17][95] = 16'sd-7;
        fc2_weights[17][96] = 16'sd23;
        fc2_weights[17][97] = 16'sd-60;
        fc2_weights[17][98] = 16'sd5;
        fc2_weights[17][99] = 16'sd-16;
        fc2_weights[17][100] = 16'sd-11;
        fc2_weights[17][101] = 16'sd-12;
        fc2_weights[17][102] = 16'sd2;
        fc2_weights[17][103] = 16'sd-36;
        fc2_weights[17][104] = 16'sd43;
        fc2_weights[17][105] = 16'sd-29;
        fc2_weights[17][106] = 16'sd-48;
        fc2_weights[17][107] = 16'sd57;
        fc2_weights[17][108] = 16'sd21;
        fc2_weights[17][109] = 16'sd-2;
        fc2_weights[17][110] = 16'sd37;
        fc2_weights[17][111] = 16'sd15;
        fc2_weights[17][112] = 16'sd-37;
        fc2_weights[17][113] = 16'sd-52;
        fc2_weights[17][114] = 16'sd-34;
        fc2_weights[17][115] = 16'sd-31;
        fc2_weights[17][116] = 16'sd42;
        fc2_weights[17][117] = 16'sd7;
        fc2_weights[17][118] = 16'sd-60;
        fc2_weights[17][119] = 16'sd4;
        fc2_weights[17][120] = 16'sd-36;
        fc2_weights[17][121] = 16'sd-11;
        fc2_weights[17][122] = 16'sd14;
        fc2_weights[17][123] = 16'sd66;
        fc2_weights[17][124] = 16'sd-51;
        fc2_weights[17][125] = 16'sd19;
        fc2_weights[17][126] = 16'sd21;
        fc2_weights[17][127] = 16'sd7;
        fc2_weights[18][0] = 16'sd-4;
        fc2_weights[18][1] = 16'sd-15;
        fc2_weights[18][2] = 16'sd15;
        fc2_weights[18][3] = 16'sd20;
        fc2_weights[18][4] = 16'sd-11;
        fc2_weights[18][5] = 16'sd13;
        fc2_weights[18][6] = 16'sd-55;
        fc2_weights[18][7] = 16'sd-26;
        fc2_weights[18][8] = 16'sd-45;
        fc2_weights[18][9] = 16'sd-17;
        fc2_weights[18][10] = 16'sd-15;
        fc2_weights[18][11] = 16'sd-23;
        fc2_weights[18][12] = 16'sd10;
        fc2_weights[18][13] = 16'sd32;
        fc2_weights[18][14] = 16'sd56;
        fc2_weights[18][15] = 16'sd36;
        fc2_weights[18][16] = 16'sd-5;
        fc2_weights[18][17] = 16'sd46;
        fc2_weights[18][18] = 16'sd-7;
        fc2_weights[18][19] = 16'sd25;
        fc2_weights[18][20] = 16'sd19;
        fc2_weights[18][21] = 16'sd-5;
        fc2_weights[18][22] = 16'sd-33;
        fc2_weights[18][23] = 16'sd11;
        fc2_weights[18][24] = 16'sd-2;
        fc2_weights[18][25] = 16'sd34;
        fc2_weights[18][26] = 16'sd-42;
        fc2_weights[18][27] = 16'sd18;
        fc2_weights[18][28] = 16'sd-24;
        fc2_weights[18][29] = 16'sd-30;
        fc2_weights[18][30] = 16'sd30;
        fc2_weights[18][31] = 16'sd-15;
        fc2_weights[18][32] = 16'sd-38;
        fc2_weights[18][33] = 16'sd-1;
        fc2_weights[18][34] = 16'sd73;
        fc2_weights[18][35] = 16'sd55;
        fc2_weights[18][36] = 16'sd-25;
        fc2_weights[18][37] = 16'sd2;
        fc2_weights[18][38] = 16'sd-23;
        fc2_weights[18][39] = 16'sd-37;
        fc2_weights[18][40] = 16'sd-4;
        fc2_weights[18][41] = 16'sd12;
        fc2_weights[18][42] = 16'sd20;
        fc2_weights[18][43] = 16'sd23;
        fc2_weights[18][44] = 16'sd48;
        fc2_weights[18][45] = 16'sd10;
        fc2_weights[18][46] = 16'sd68;
        fc2_weights[18][47] = 16'sd-16;
        fc2_weights[18][48] = 16'sd59;
        fc2_weights[18][49] = 16'sd4;
        fc2_weights[18][50] = 16'sd73;
        fc2_weights[18][51] = 16'sd-7;
        fc2_weights[18][52] = 16'sd76;
        fc2_weights[18][53] = 16'sd-31;
        fc2_weights[18][54] = 16'sd-26;
        fc2_weights[18][55] = 16'sd-19;
        fc2_weights[18][56] = 16'sd6;
        fc2_weights[18][57] = 16'sd16;
        fc2_weights[18][58] = 16'sd30;
        fc2_weights[18][59] = 16'sd22;
        fc2_weights[18][60] = 16'sd1;
        fc2_weights[18][61] = 16'sd-51;
        fc2_weights[18][62] = 16'sd34;
        fc2_weights[18][63] = 16'sd29;
        fc2_weights[18][64] = 16'sd-44;
        fc2_weights[18][65] = 16'sd40;
        fc2_weights[18][66] = 16'sd-12;
        fc2_weights[18][67] = 16'sd-10;
        fc2_weights[18][68] = 16'sd36;
        fc2_weights[18][69] = 16'sd17;
        fc2_weights[18][70] = 16'sd-14;
        fc2_weights[18][71] = 16'sd27;
        fc2_weights[18][72] = 16'sd25;
        fc2_weights[18][73] = 16'sd-34;
        fc2_weights[18][74] = 16'sd36;
        fc2_weights[18][75] = 16'sd11;
        fc2_weights[18][76] = 16'sd-35;
        fc2_weights[18][77] = 16'sd15;
        fc2_weights[18][78] = 16'sd35;
        fc2_weights[18][79] = 16'sd-7;
        fc2_weights[18][80] = 16'sd-30;
        fc2_weights[18][81] = 16'sd7;
        fc2_weights[18][82] = 16'sd-24;
        fc2_weights[18][83] = 16'sd-24;
        fc2_weights[18][84] = 16'sd38;
        fc2_weights[18][85] = 16'sd-19;
        fc2_weights[18][86] = 16'sd-7;
        fc2_weights[18][87] = 16'sd-20;
        fc2_weights[18][88] = 16'sd42;
        fc2_weights[18][89] = 16'sd-41;
        fc2_weights[18][90] = 16'sd44;
        fc2_weights[18][91] = 16'sd23;
        fc2_weights[18][92] = 16'sd36;
        fc2_weights[18][93] = 16'sd-42;
        fc2_weights[18][94] = 16'sd27;
        fc2_weights[18][95] = 16'sd-23;
        fc2_weights[18][96] = 16'sd39;
        fc2_weights[18][97] = 16'sd-4;
        fc2_weights[18][98] = 16'sd-45;
        fc2_weights[18][99] = 16'sd-19;
        fc2_weights[18][100] = 16'sd0;
        fc2_weights[18][101] = 16'sd11;
        fc2_weights[18][102] = 16'sd31;
        fc2_weights[18][103] = 16'sd12;
        fc2_weights[18][104] = 16'sd42;
        fc2_weights[18][105] = 16'sd-11;
        fc2_weights[18][106] = 16'sd3;
        fc2_weights[18][107] = 16'sd38;
        fc2_weights[18][108] = 16'sd-17;
        fc2_weights[18][109] = 16'sd-45;
        fc2_weights[18][110] = 16'sd27;
        fc2_weights[18][111] = 16'sd-21;
        fc2_weights[18][112] = 16'sd-36;
        fc2_weights[18][113] = 16'sd-30;
        fc2_weights[18][114] = 16'sd-16;
        fc2_weights[18][115] = 16'sd-53;
        fc2_weights[18][116] = 16'sd-18;
        fc2_weights[18][117] = 16'sd-32;
        fc2_weights[18][118] = 16'sd-23;
        fc2_weights[18][119] = 16'sd-12;
        fc2_weights[18][120] = 16'sd-26;
        fc2_weights[18][121] = 16'sd1;
        fc2_weights[18][122] = 16'sd43;
        fc2_weights[18][123] = 16'sd38;
        fc2_weights[18][124] = 16'sd-22;
        fc2_weights[18][125] = 16'sd31;
        fc2_weights[18][126] = 16'sd41;
        fc2_weights[18][127] = 16'sd-18;
        fc2_weights[19][0] = 16'sd-16;
        fc2_weights[19][1] = 16'sd-44;
        fc2_weights[19][2] = 16'sd-29;
        fc2_weights[19][3] = 16'sd34;
        fc2_weights[19][4] = 16'sd-38;
        fc2_weights[19][5] = 16'sd9;
        fc2_weights[19][6] = 16'sd-47;
        fc2_weights[19][7] = 16'sd-29;
        fc2_weights[19][8] = 16'sd-40;
        fc2_weights[19][9] = 16'sd25;
        fc2_weights[19][10] = 16'sd-17;
        fc2_weights[19][11] = 16'sd-12;
        fc2_weights[19][12] = 16'sd-27;
        fc2_weights[19][13] = 16'sd4;
        fc2_weights[19][14] = 16'sd15;
        fc2_weights[19][15] = 16'sd33;
        fc2_weights[19][16] = 16'sd16;
        fc2_weights[19][17] = 16'sd36;
        fc2_weights[19][18] = 16'sd-15;
        fc2_weights[19][19] = 16'sd-22;
        fc2_weights[19][20] = 16'sd2;
        fc2_weights[19][21] = 16'sd-61;
        fc2_weights[19][22] = 16'sd-26;
        fc2_weights[19][23] = 16'sd-15;
        fc2_weights[19][24] = 16'sd8;
        fc2_weights[19][25] = 16'sd-12;
        fc2_weights[19][26] = 16'sd4;
        fc2_weights[19][27] = 16'sd25;
        fc2_weights[19][28] = 16'sd1;
        fc2_weights[19][29] = 16'sd-29;
        fc2_weights[19][30] = 16'sd6;
        fc2_weights[19][31] = 16'sd-20;
        fc2_weights[19][32] = 16'sd-17;
        fc2_weights[19][33] = 16'sd-43;
        fc2_weights[19][34] = 16'sd25;
        fc2_weights[19][35] = 16'sd63;
        fc2_weights[19][36] = 16'sd-44;
        fc2_weights[19][37] = 16'sd-13;
        fc2_weights[19][38] = 16'sd-3;
        fc2_weights[19][39] = 16'sd-47;
        fc2_weights[19][40] = 16'sd-6;
        fc2_weights[19][41] = 16'sd3;
        fc2_weights[19][42] = 16'sd-23;
        fc2_weights[19][43] = 16'sd0;
        fc2_weights[19][44] = 16'sd35;
        fc2_weights[19][45] = 16'sd20;
        fc2_weights[19][46] = 16'sd-38;
        fc2_weights[19][47] = 16'sd12;
        fc2_weights[19][48] = 16'sd-7;
        fc2_weights[19][49] = 16'sd-18;
        fc2_weights[19][50] = 16'sd32;
        fc2_weights[19][51] = 16'sd21;
        fc2_weights[19][52] = 16'sd21;
        fc2_weights[19][53] = 16'sd-51;
        fc2_weights[19][54] = 16'sd-55;
        fc2_weights[19][55] = 16'sd5;
        fc2_weights[19][56] = 16'sd18;
        fc2_weights[19][57] = 16'sd34;
        fc2_weights[19][58] = 16'sd12;
        fc2_weights[19][59] = 16'sd4;
        fc2_weights[19][60] = 16'sd11;
        fc2_weights[19][61] = 16'sd-35;
        fc2_weights[19][62] = 16'sd7;
        fc2_weights[19][63] = 16'sd0;
        fc2_weights[19][64] = 16'sd-53;
        fc2_weights[19][65] = 16'sd33;
        fc2_weights[19][66] = 16'sd31;
        fc2_weights[19][67] = 16'sd-34;
        fc2_weights[19][68] = 16'sd22;
        fc2_weights[19][69] = 16'sd60;
        fc2_weights[19][70] = 16'sd-38;
        fc2_weights[19][71] = 16'sd-42;
        fc2_weights[19][72] = 16'sd-65;
        fc2_weights[19][73] = 16'sd-25;
        fc2_weights[19][74] = 16'sd21;
        fc2_weights[19][75] = 16'sd-8;
        fc2_weights[19][76] = 16'sd11;
        fc2_weights[19][77] = 16'sd21;
        fc2_weights[19][78] = 16'sd25;
        fc2_weights[19][79] = 16'sd-26;
        fc2_weights[19][80] = 16'sd-55;
        fc2_weights[19][81] = 16'sd19;
        fc2_weights[19][82] = 16'sd-51;
        fc2_weights[19][83] = 16'sd-50;
        fc2_weights[19][84] = 16'sd-32;
        fc2_weights[19][85] = 16'sd-5;
        fc2_weights[19][86] = 16'sd-26;
        fc2_weights[19][87] = 16'sd-39;
        fc2_weights[19][88] = 16'sd2;
        fc2_weights[19][89] = 16'sd-64;
        fc2_weights[19][90] = 16'sd-4;
        fc2_weights[19][91] = 16'sd8;
        fc2_weights[19][92] = 16'sd3;
        fc2_weights[19][93] = 16'sd-13;
        fc2_weights[19][94] = 16'sd27;
        fc2_weights[19][95] = 16'sd-32;
        fc2_weights[19][96] = 16'sd38;
        fc2_weights[19][97] = 16'sd-29;
        fc2_weights[19][98] = 16'sd-14;
        fc2_weights[19][99] = 16'sd-30;
        fc2_weights[19][100] = 16'sd15;
        fc2_weights[19][101] = 16'sd-3;
        fc2_weights[19][102] = 16'sd-11;
        fc2_weights[19][103] = 16'sd-24;
        fc2_weights[19][104] = 16'sd11;
        fc2_weights[19][105] = 16'sd-36;
        fc2_weights[19][106] = 16'sd-17;
        fc2_weights[19][107] = 16'sd32;
        fc2_weights[19][108] = 16'sd-33;
        fc2_weights[19][109] = 16'sd-18;
        fc2_weights[19][110] = 16'sd33;
        fc2_weights[19][111] = 16'sd-25;
        fc2_weights[19][112] = 16'sd-18;
        fc2_weights[19][113] = 16'sd-57;
        fc2_weights[19][114] = 16'sd0;
        fc2_weights[19][115] = 16'sd-26;
        fc2_weights[19][116] = 16'sd-23;
        fc2_weights[19][117] = 16'sd-9;
        fc2_weights[19][118] = 16'sd-60;
        fc2_weights[19][119] = 16'sd23;
        fc2_weights[19][120] = 16'sd-51;
        fc2_weights[19][121] = 16'sd-43;
        fc2_weights[19][122] = 16'sd6;
        fc2_weights[19][123] = 16'sd39;
        fc2_weights[19][124] = 16'sd-27;
        fc2_weights[19][125] = 16'sd20;
        fc2_weights[19][126] = 16'sd16;
        fc2_weights[19][127] = 16'sd-51;
        fc2_weights[20][0] = 16'sd-73;
        fc2_weights[20][1] = 16'sd-19;
        fc2_weights[20][2] = 16'sd61;
        fc2_weights[20][3] = 16'sd-11;
        fc2_weights[20][4] = 16'sd-62;
        fc2_weights[20][5] = 16'sd-107;
        fc2_weights[20][6] = 16'sd-40;
        fc2_weights[20][7] = 16'sd29;
        fc2_weights[20][8] = 16'sd-69;
        fc2_weights[20][9] = 16'sd-23;
        fc2_weights[20][10] = 16'sd-20;
        fc2_weights[20][11] = 16'sd-59;
        fc2_weights[20][12] = 16'sd-27;
        fc2_weights[20][13] = 16'sd-59;
        fc2_weights[20][14] = 16'sd20;
        fc2_weights[20][15] = 16'sd36;
        fc2_weights[20][16] = 16'sd27;
        fc2_weights[20][17] = 16'sd-5;
        fc2_weights[20][18] = 16'sd-17;
        fc2_weights[20][19] = 16'sd9;
        fc2_weights[20][20] = 16'sd17;
        fc2_weights[20][21] = 16'sd15;
        fc2_weights[20][22] = 16'sd-5;
        fc2_weights[20][23] = 16'sd-35;
        fc2_weights[20][24] = 16'sd60;
        fc2_weights[20][25] = 16'sd-10;
        fc2_weights[20][26] = 16'sd11;
        fc2_weights[20][27] = 16'sd-11;
        fc2_weights[20][28] = 16'sd-34;
        fc2_weights[20][29] = 16'sd-13;
        fc2_weights[20][30] = 16'sd-26;
        fc2_weights[20][31] = 16'sd-65;
        fc2_weights[20][32] = 16'sd40;
        fc2_weights[20][33] = 16'sd-47;
        fc2_weights[20][34] = 16'sd32;
        fc2_weights[20][35] = 16'sd9;
        fc2_weights[20][36] = 16'sd-8;
        fc2_weights[20][37] = 16'sd23;
        fc2_weights[20][38] = 16'sd-52;
        fc2_weights[20][39] = 16'sd-59;
        fc2_weights[20][40] = 16'sd-12;
        fc2_weights[20][41] = 16'sd11;
        fc2_weights[20][42] = 16'sd-57;
        fc2_weights[20][43] = 16'sd10;
        fc2_weights[20][44] = 16'sd40;
        fc2_weights[20][45] = 16'sd100;
        fc2_weights[20][46] = 16'sd18;
        fc2_weights[20][47] = 16'sd4;
        fc2_weights[20][48] = 16'sd-16;
        fc2_weights[20][49] = 16'sd-7;
        fc2_weights[20][50] = 16'sd49;
        fc2_weights[20][51] = 16'sd-72;
        fc2_weights[20][52] = 16'sd29;
        fc2_weights[20][53] = 16'sd-16;
        fc2_weights[20][54] = 16'sd-26;
        fc2_weights[20][55] = 16'sd1;
        fc2_weights[20][56] = 16'sd23;
        fc2_weights[20][57] = 16'sd69;
        fc2_weights[20][58] = 16'sd34;
        fc2_weights[20][59] = 16'sd64;
        fc2_weights[20][60] = 16'sd-8;
        fc2_weights[20][61] = 16'sd9;
        fc2_weights[20][62] = 16'sd41;
        fc2_weights[20][63] = 16'sd41;
        fc2_weights[20][64] = 16'sd-20;
        fc2_weights[20][65] = 16'sd37;
        fc2_weights[20][66] = 16'sd47;
        fc2_weights[20][67] = 16'sd-37;
        fc2_weights[20][68] = 16'sd-22;
        fc2_weights[20][69] = 16'sd94;
        fc2_weights[20][70] = 16'sd-41;
        fc2_weights[20][71] = 16'sd4;
        fc2_weights[20][72] = 16'sd-34;
        fc2_weights[20][73] = 16'sd-50;
        fc2_weights[20][74] = 16'sd17;
        fc2_weights[20][75] = 16'sd-14;
        fc2_weights[20][76] = 16'sd-34;
        fc2_weights[20][77] = 16'sd-23;
        fc2_weights[20][78] = 16'sd-20;
        fc2_weights[20][79] = 16'sd-9;
        fc2_weights[20][80] = 16'sd-43;
        fc2_weights[20][81] = 16'sd-2;
        fc2_weights[20][82] = 16'sd-24;
        fc2_weights[20][83] = 16'sd21;
        fc2_weights[20][84] = 16'sd5;
        fc2_weights[20][85] = 16'sd-34;
        fc2_weights[20][86] = 16'sd-12;
        fc2_weights[20][87] = 16'sd-34;
        fc2_weights[20][88] = 16'sd79;
        fc2_weights[20][89] = 16'sd-56;
        fc2_weights[20][90] = 16'sd43;
        fc2_weights[20][91] = 16'sd25;
        fc2_weights[20][92] = 16'sd10;
        fc2_weights[20][93] = 16'sd-70;
        fc2_weights[20][94] = 16'sd-48;
        fc2_weights[20][95] = 16'sd12;
        fc2_weights[20][96] = 16'sd51;
        fc2_weights[20][97] = 16'sd-19;
        fc2_weights[20][98] = 16'sd-2;
        fc2_weights[20][99] = 16'sd-28;
        fc2_weights[20][100] = 16'sd-10;
        fc2_weights[20][101] = 16'sd-3;
        fc2_weights[20][102] = 16'sd31;
        fc2_weights[20][103] = 16'sd-18;
        fc2_weights[20][104] = 16'sd24;
        fc2_weights[20][105] = 16'sd-33;
        fc2_weights[20][106] = 16'sd-34;
        fc2_weights[20][107] = 16'sd25;
        fc2_weights[20][108] = 16'sd-53;
        fc2_weights[20][109] = 16'sd-45;
        fc2_weights[20][110] = 16'sd27;
        fc2_weights[20][111] = 16'sd16;
        fc2_weights[20][112] = 16'sd-67;
        fc2_weights[20][113] = 16'sd-81;
        fc2_weights[20][114] = 16'sd-39;
        fc2_weights[20][115] = 16'sd-35;
        fc2_weights[20][116] = 16'sd65;
        fc2_weights[20][117] = 16'sd62;
        fc2_weights[20][118] = 16'sd-62;
        fc2_weights[20][119] = 16'sd-23;
        fc2_weights[20][120] = 16'sd-3;
        fc2_weights[20][121] = 16'sd-6;
        fc2_weights[20][122] = 16'sd-5;
        fc2_weights[20][123] = 16'sd48;
        fc2_weights[20][124] = 16'sd-6;
        fc2_weights[20][125] = 16'sd37;
        fc2_weights[20][126] = 16'sd36;
        fc2_weights[20][127] = 16'sd5;
        fc2_weights[21][0] = 16'sd1;
        fc2_weights[21][1] = 16'sd-94;
        fc2_weights[21][2] = 16'sd8;
        fc2_weights[21][3] = 16'sd-27;
        fc2_weights[21][4] = 16'sd-17;
        fc2_weights[21][5] = 16'sd17;
        fc2_weights[21][6] = 16'sd-14;
        fc2_weights[21][7] = 16'sd-30;
        fc2_weights[21][8] = 16'sd71;
        fc2_weights[21][9] = 16'sd-5;
        fc2_weights[21][10] = 16'sd-10;
        fc2_weights[21][11] = 16'sd-100;
        fc2_weights[21][12] = 16'sd-35;
        fc2_weights[21][13] = 16'sd16;
        fc2_weights[21][14] = 16'sd80;
        fc2_weights[21][15] = 16'sd-7;
        fc2_weights[21][16] = 16'sd-28;
        fc2_weights[21][17] = 16'sd11;
        fc2_weights[21][18] = 16'sd55;
        fc2_weights[21][19] = 16'sd2;
        fc2_weights[21][20] = 16'sd0;
        fc2_weights[21][21] = 16'sd-25;
        fc2_weights[21][22] = 16'sd-6;
        fc2_weights[21][23] = 16'sd-22;
        fc2_weights[21][24] = 16'sd-4;
        fc2_weights[21][25] = 16'sd70;
        fc2_weights[21][26] = 16'sd-74;
        fc2_weights[21][27] = 16'sd18;
        fc2_weights[21][28] = 16'sd-29;
        fc2_weights[21][29] = 16'sd-45;
        fc2_weights[21][30] = 16'sd3;
        fc2_weights[21][31] = 16'sd-50;
        fc2_weights[21][32] = 16'sd-41;
        fc2_weights[21][33] = 16'sd-31;
        fc2_weights[21][34] = 16'sd19;
        fc2_weights[21][35] = 16'sd-17;
        fc2_weights[21][36] = 16'sd-37;
        fc2_weights[21][37] = 16'sd17;
        fc2_weights[21][38] = 16'sd-40;
        fc2_weights[21][39] = 16'sd-48;
        fc2_weights[21][40] = 16'sd-32;
        fc2_weights[21][41] = 16'sd83;
        fc2_weights[21][42] = 16'sd-6;
        fc2_weights[21][43] = 16'sd29;
        fc2_weights[21][44] = 16'sd2;
        fc2_weights[21][45] = 16'sd10;
        fc2_weights[21][46] = 16'sd4;
        fc2_weights[21][47] = 16'sd-40;
        fc2_weights[21][48] = 16'sd111;
        fc2_weights[21][49] = 16'sd-2;
        fc2_weights[21][50] = 16'sd47;
        fc2_weights[21][51] = 16'sd-11;
        fc2_weights[21][52] = 16'sd20;
        fc2_weights[21][53] = 16'sd10;
        fc2_weights[21][54] = 16'sd43;
        fc2_weights[21][55] = 16'sd56;
        fc2_weights[21][56] = 16'sd-6;
        fc2_weights[21][57] = 16'sd-33;
        fc2_weights[21][58] = 16'sd39;
        fc2_weights[21][59] = 16'sd43;
        fc2_weights[21][60] = 16'sd8;
        fc2_weights[21][61] = 16'sd-74;
        fc2_weights[21][62] = 16'sd-18;
        fc2_weights[21][63] = 16'sd38;
        fc2_weights[21][64] = 16'sd-5;
        fc2_weights[21][65] = 16'sd45;
        fc2_weights[21][66] = 16'sd-5;
        fc2_weights[21][67] = 16'sd-19;
        fc2_weights[21][68] = 16'sd-1;
        fc2_weights[21][69] = 16'sd35;
        fc2_weights[21][70] = 16'sd11;
        fc2_weights[21][71] = 16'sd-10;
        fc2_weights[21][72] = 16'sd65;
        fc2_weights[21][73] = 16'sd-9;
        fc2_weights[21][74] = 16'sd16;
        fc2_weights[21][75] = 16'sd-23;
        fc2_weights[21][76] = 16'sd-23;
        fc2_weights[21][77] = 16'sd-14;
        fc2_weights[21][78] = 16'sd1;
        fc2_weights[21][79] = 16'sd-30;
        fc2_weights[21][80] = 16'sd-16;
        fc2_weights[21][81] = 16'sd68;
        fc2_weights[21][82] = 16'sd-14;
        fc2_weights[21][83] = 16'sd-8;
        fc2_weights[21][84] = 16'sd31;
        fc2_weights[21][85] = 16'sd14;
        fc2_weights[21][86] = 16'sd-26;
        fc2_weights[21][87] = 16'sd-93;
        fc2_weights[21][88] = 16'sd60;
        fc2_weights[21][89] = 16'sd-31;
        fc2_weights[21][90] = 16'sd1;
        fc2_weights[21][91] = 16'sd20;
        fc2_weights[21][92] = 16'sd17;
        fc2_weights[21][93] = 16'sd-63;
        fc2_weights[21][94] = 16'sd35;
        fc2_weights[21][95] = 16'sd-14;
        fc2_weights[21][96] = 16'sd11;
        fc2_weights[21][97] = 16'sd8;
        fc2_weights[21][98] = 16'sd23;
        fc2_weights[21][99] = 16'sd10;
        fc2_weights[21][100] = 16'sd27;
        fc2_weights[21][101] = 16'sd-32;
        fc2_weights[21][102] = 16'sd24;
        fc2_weights[21][103] = 16'sd58;
        fc2_weights[21][104] = 16'sd-13;
        fc2_weights[21][105] = 16'sd30;
        fc2_weights[21][106] = 16'sd6;
        fc2_weights[21][107] = 16'sd41;
        fc2_weights[21][108] = 16'sd15;
        fc2_weights[21][109] = 16'sd-47;
        fc2_weights[21][110] = 16'sd70;
        fc2_weights[21][111] = 16'sd-11;
        fc2_weights[21][112] = 16'sd38;
        fc2_weights[21][113] = 16'sd-57;
        fc2_weights[21][114] = 16'sd38;
        fc2_weights[21][115] = 16'sd-14;
        fc2_weights[21][116] = 16'sd27;
        fc2_weights[21][117] = 16'sd42;
        fc2_weights[21][118] = 16'sd-40;
        fc2_weights[21][119] = 16'sd-1;
        fc2_weights[21][120] = 16'sd19;
        fc2_weights[21][121] = 16'sd33;
        fc2_weights[21][122] = 16'sd103;
        fc2_weights[21][123] = 16'sd28;
        fc2_weights[21][124] = 16'sd-8;
        fc2_weights[21][125] = 16'sd19;
        fc2_weights[21][126] = 16'sd38;
        fc2_weights[21][127] = 16'sd-5;
        fc2_weights[22][0] = 16'sd41;
        fc2_weights[22][1] = 16'sd25;
        fc2_weights[22][2] = 16'sd-8;
        fc2_weights[22][3] = 16'sd-41;
        fc2_weights[22][4] = 16'sd25;
        fc2_weights[22][5] = 16'sd15;
        fc2_weights[22][6] = 16'sd25;
        fc2_weights[22][7] = 16'sd42;
        fc2_weights[22][8] = 16'sd25;
        fc2_weights[22][9] = 16'sd39;
        fc2_weights[22][10] = 16'sd-27;
        fc2_weights[22][11] = 16'sd-24;
        fc2_weights[22][12] = 16'sd-7;
        fc2_weights[22][13] = 16'sd-42;
        fc2_weights[22][14] = 16'sd29;
        fc2_weights[22][15] = 16'sd-46;
        fc2_weights[22][16] = 16'sd-6;
        fc2_weights[22][17] = 16'sd-42;
        fc2_weights[22][18] = 16'sd48;
        fc2_weights[22][19] = 16'sd-6;
        fc2_weights[22][20] = 16'sd-57;
        fc2_weights[22][21] = 16'sd-36;
        fc2_weights[22][22] = 16'sd66;
        fc2_weights[22][23] = 16'sd38;
        fc2_weights[22][24] = 16'sd3;
        fc2_weights[22][25] = 16'sd-26;
        fc2_weights[22][26] = 16'sd-27;
        fc2_weights[22][27] = 16'sd26;
        fc2_weights[22][28] = 16'sd-20;
        fc2_weights[22][29] = 16'sd39;
        fc2_weights[22][30] = 16'sd-13;
        fc2_weights[22][31] = 16'sd18;
        fc2_weights[22][32] = 16'sd-9;
        fc2_weights[22][33] = 16'sd-14;
        fc2_weights[22][34] = 16'sd-51;
        fc2_weights[22][35] = 16'sd-4;
        fc2_weights[22][36] = 16'sd91;
        fc2_weights[22][37] = 16'sd-8;
        fc2_weights[22][38] = 16'sd39;
        fc2_weights[22][39] = 16'sd22;
        fc2_weights[22][40] = 16'sd-44;
        fc2_weights[22][41] = 16'sd8;
        fc2_weights[22][42] = 16'sd2;
        fc2_weights[22][43] = 16'sd2;
        fc2_weights[22][44] = 16'sd-50;
        fc2_weights[22][45] = 16'sd-23;
        fc2_weights[22][46] = 16'sd38;
        fc2_weights[22][47] = 16'sd37;
        fc2_weights[22][48] = 16'sd5;
        fc2_weights[22][49] = 16'sd53;
        fc2_weights[22][50] = 16'sd8;
        fc2_weights[22][51] = 16'sd-1;
        fc2_weights[22][52] = 16'sd-11;
        fc2_weights[22][53] = 16'sd-10;
        fc2_weights[22][54] = 16'sd-22;
        fc2_weights[22][55] = 16'sd-14;
        fc2_weights[22][56] = 16'sd4;
        fc2_weights[22][57] = 16'sd-53;
        fc2_weights[22][58] = 16'sd-43;
        fc2_weights[22][59] = 16'sd-73;
        fc2_weights[22][60] = 16'sd21;
        fc2_weights[22][61] = 16'sd-9;
        fc2_weights[22][62] = 16'sd55;
        fc2_weights[22][63] = 16'sd-25;
        fc2_weights[22][64] = 16'sd23;
        fc2_weights[22][65] = 16'sd1;
        fc2_weights[22][66] = 16'sd-10;
        fc2_weights[22][67] = 16'sd46;
        fc2_weights[22][68] = 16'sd-42;
        fc2_weights[22][69] = 16'sd-79;
        fc2_weights[22][70] = 16'sd8;
        fc2_weights[22][71] = 16'sd-66;
        fc2_weights[22][72] = 16'sd17;
        fc2_weights[22][73] = 16'sd23;
        fc2_weights[22][74] = 16'sd8;
        fc2_weights[22][75] = 16'sd13;
        fc2_weights[22][76] = 16'sd-17;
        fc2_weights[22][77] = 16'sd95;
        fc2_weights[22][78] = 16'sd-29;
        fc2_weights[22][79] = 16'sd15;
        fc2_weights[22][80] = 16'sd-38;
        fc2_weights[22][81] = 16'sd39;
        fc2_weights[22][82] = 16'sd44;
        fc2_weights[22][83] = 16'sd-67;
        fc2_weights[22][84] = 16'sd-33;
        fc2_weights[22][85] = 16'sd37;
        fc2_weights[22][86] = 16'sd44;
        fc2_weights[22][87] = 16'sd-30;
        fc2_weights[22][88] = 16'sd9;
        fc2_weights[22][89] = 16'sd46;
        fc2_weights[22][90] = 16'sd-51;
        fc2_weights[22][91] = 16'sd11;
        fc2_weights[22][92] = 16'sd110;
        fc2_weights[22][93] = 16'sd32;
        fc2_weights[22][94] = 16'sd-39;
        fc2_weights[22][95] = 16'sd-52;
        fc2_weights[22][96] = 16'sd-75;
        fc2_weights[22][97] = 16'sd78;
        fc2_weights[22][98] = 16'sd31;
        fc2_weights[22][99] = 16'sd49;
        fc2_weights[22][100] = 16'sd-28;
        fc2_weights[22][101] = 16'sd18;
        fc2_weights[22][102] = 16'sd-35;
        fc2_weights[22][103] = 16'sd-67;
        fc2_weights[22][104] = 16'sd-6;
        fc2_weights[22][105] = 16'sd9;
        fc2_weights[22][106] = 16'sd31;
        fc2_weights[22][107] = 16'sd13;
        fc2_weights[22][108] = 16'sd73;
        fc2_weights[22][109] = 16'sd25;
        fc2_weights[22][110] = 16'sd-33;
        fc2_weights[22][111] = 16'sd31;
        fc2_weights[22][112] = 16'sd8;
        fc2_weights[22][113] = 16'sd55;
        fc2_weights[22][114] = 16'sd17;
        fc2_weights[22][115] = 16'sd54;
        fc2_weights[22][116] = 16'sd-14;
        fc2_weights[22][117] = 16'sd-16;
        fc2_weights[22][118] = 16'sd59;
        fc2_weights[22][119] = 16'sd-59;
        fc2_weights[22][120] = 16'sd-29;
        fc2_weights[22][121] = 16'sd3;
        fc2_weights[22][122] = 16'sd-22;
        fc2_weights[22][123] = 16'sd15;
        fc2_weights[22][124] = 16'sd-18;
        fc2_weights[22][125] = 16'sd-47;
        fc2_weights[22][126] = 16'sd-10;
        fc2_weights[22][127] = 16'sd-13;
        fc2_weights[23][0] = 16'sd26;
        fc2_weights[23][1] = 16'sd25;
        fc2_weights[23][2] = 16'sd-32;
        fc2_weights[23][3] = 16'sd119;
        fc2_weights[23][4] = 16'sd-14;
        fc2_weights[23][5] = 16'sd-7;
        fc2_weights[23][6] = 16'sd19;
        fc2_weights[23][7] = 16'sd-21;
        fc2_weights[23][8] = 16'sd56;
        fc2_weights[23][9] = 16'sd39;
        fc2_weights[23][10] = 16'sd7;
        fc2_weights[23][11] = 16'sd-3;
        fc2_weights[23][12] = 16'sd66;
        fc2_weights[23][13] = 16'sd-7;
        fc2_weights[23][14] = 16'sd-87;
        fc2_weights[23][15] = 16'sd-2;
        fc2_weights[23][16] = 16'sd-41;
        fc2_weights[23][17] = 16'sd30;
        fc2_weights[23][18] = 16'sd2;
        fc2_weights[23][19] = 16'sd-8;
        fc2_weights[23][20] = 16'sd10;
        fc2_weights[23][21] = 16'sd-36;
        fc2_weights[23][22] = 16'sd19;
        fc2_weights[23][23] = 16'sd-76;
        fc2_weights[23][24] = 16'sd-25;
        fc2_weights[23][25] = 16'sd-74;
        fc2_weights[23][26] = 16'sd-11;
        fc2_weights[23][27] = 16'sd-34;
        fc2_weights[23][28] = 16'sd74;
        fc2_weights[23][29] = 16'sd11;
        fc2_weights[23][30] = 16'sd26;
        fc2_weights[23][31] = 16'sd-23;
        fc2_weights[23][32] = 16'sd62;
        fc2_weights[23][33] = 16'sd46;
        fc2_weights[23][34] = 16'sd13;
        fc2_weights[23][35] = 16'sd-53;
        fc2_weights[23][36] = 16'sd49;
        fc2_weights[23][37] = 16'sd17;
        fc2_weights[23][38] = 16'sd-27;
        fc2_weights[23][39] = 16'sd46;
        fc2_weights[23][40] = 16'sd-45;
        fc2_weights[23][41] = 16'sd-76;
        fc2_weights[23][42] = 16'sd-33;
        fc2_weights[23][43] = 16'sd21;
        fc2_weights[23][44] = 16'sd-39;
        fc2_weights[23][45] = 16'sd-50;
        fc2_weights[23][46] = 16'sd-49;
        fc2_weights[23][47] = 16'sd12;
        fc2_weights[23][48] = 16'sd-1;
        fc2_weights[23][49] = 16'sd-10;
        fc2_weights[23][50] = 16'sd-41;
        fc2_weights[23][51] = 16'sd-26;
        fc2_weights[23][52] = 16'sd42;
        fc2_weights[23][53] = 16'sd26;
        fc2_weights[23][54] = 16'sd-17;
        fc2_weights[23][55] = 16'sd23;
        fc2_weights[23][56] = 16'sd-14;
        fc2_weights[23][57] = 16'sd-64;
        fc2_weights[23][58] = 16'sd-78;
        fc2_weights[23][59] = 16'sd18;
        fc2_weights[23][60] = 16'sd-17;
        fc2_weights[23][61] = 16'sd23;
        fc2_weights[23][62] = 16'sd-78;
        fc2_weights[23][63] = 16'sd2;
        fc2_weights[23][64] = 16'sd-2;
        fc2_weights[23][65] = 16'sd-40;
        fc2_weights[23][66] = 16'sd-13;
        fc2_weights[23][67] = 16'sd-33;
        fc2_weights[23][68] = 16'sd11;
        fc2_weights[23][69] = 16'sd-26;
        fc2_weights[23][70] = 16'sd-10;
        fc2_weights[23][71] = 16'sd-39;
        fc2_weights[23][72] = 16'sd5;
        fc2_weights[23][73] = 16'sd34;
        fc2_weights[23][74] = 16'sd21;
        fc2_weights[23][75] = 16'sd-30;
        fc2_weights[23][76] = 16'sd11;
        fc2_weights[23][77] = 16'sd-18;
        fc2_weights[23][78] = 16'sd-31;
        fc2_weights[23][79] = 16'sd-22;
        fc2_weights[23][80] = 16'sd44;
        fc2_weights[23][81] = 16'sd-61;
        fc2_weights[23][82] = 16'sd-7;
        fc2_weights[23][83] = 16'sd13;
        fc2_weights[23][84] = 16'sd-14;
        fc2_weights[23][85] = 16'sd4;
        fc2_weights[23][86] = 16'sd-24;
        fc2_weights[23][87] = 16'sd1;
        fc2_weights[23][88] = 16'sd-57;
        fc2_weights[23][89] = 16'sd-7;
        fc2_weights[23][90] = 16'sd-22;
        fc2_weights[23][91] = 16'sd-21;
        fc2_weights[23][92] = 16'sd-48;
        fc2_weights[23][93] = 16'sd47;
        fc2_weights[23][94] = 16'sd17;
        fc2_weights[23][95] = 16'sd-10;
        fc2_weights[23][96] = 16'sd-23;
        fc2_weights[23][97] = 16'sd14;
        fc2_weights[23][98] = 16'sd-37;
        fc2_weights[23][99] = 16'sd-21;
        fc2_weights[23][100] = 16'sd-98;
        fc2_weights[23][101] = 16'sd19;
        fc2_weights[23][102] = 16'sd-93;
        fc2_weights[23][103] = 16'sd-88;
        fc2_weights[23][104] = 16'sd-72;
        fc2_weights[23][105] = 16'sd-19;
        fc2_weights[23][106] = 16'sd-8;
        fc2_weights[23][107] = 16'sd-61;
        fc2_weights[23][108] = 16'sd45;
        fc2_weights[23][109] = 16'sd19;
        fc2_weights[23][110] = 16'sd-72;
        fc2_weights[23][111] = 16'sd-44;
        fc2_weights[23][112] = 16'sd4;
        fc2_weights[23][113] = 16'sd25;
        fc2_weights[23][114] = 16'sd-55;
        fc2_weights[23][115] = 16'sd15;
        fc2_weights[23][116] = 16'sd-5;
        fc2_weights[23][117] = 16'sd-10;
        fc2_weights[23][118] = 16'sd0;
        fc2_weights[23][119] = 16'sd2;
        fc2_weights[23][120] = 16'sd18;
        fc2_weights[23][121] = 16'sd-64;
        fc2_weights[23][122] = 16'sd-102;
        fc2_weights[23][123] = 16'sd-67;
        fc2_weights[23][124] = 16'sd-30;
        fc2_weights[23][125] = 16'sd-75;
        fc2_weights[23][126] = 16'sd-31;
        fc2_weights[23][127] = 16'sd-66;
        fc2_weights[24][0] = 16'sd-24;
        fc2_weights[24][1] = 16'sd-62;
        fc2_weights[24][2] = 16'sd-42;
        fc2_weights[24][3] = 16'sd-66;
        fc2_weights[24][4] = 16'sd38;
        fc2_weights[24][5] = 16'sd39;
        fc2_weights[24][6] = 16'sd39;
        fc2_weights[24][7] = 16'sd46;
        fc2_weights[24][8] = 16'sd60;
        fc2_weights[24][9] = 16'sd15;
        fc2_weights[24][10] = 16'sd-54;
        fc2_weights[24][11] = 16'sd16;
        fc2_weights[24][12] = 16'sd7;
        fc2_weights[24][13] = 16'sd-1;
        fc2_weights[24][14] = 16'sd28;
        fc2_weights[24][15] = 16'sd-23;
        fc2_weights[24][16] = 16'sd-10;
        fc2_weights[24][17] = 16'sd-26;
        fc2_weights[24][18] = 16'sd36;
        fc2_weights[24][19] = 16'sd-58;
        fc2_weights[24][20] = 16'sd-5;
        fc2_weights[24][21] = 16'sd-41;
        fc2_weights[24][22] = 16'sd60;
        fc2_weights[24][23] = 16'sd36;
        fc2_weights[24][24] = 16'sd0;
        fc2_weights[24][25] = 16'sd58;
        fc2_weights[24][26] = 16'sd-48;
        fc2_weights[24][27] = 16'sd39;
        fc2_weights[24][28] = 16'sd-7;
        fc2_weights[24][29] = 16'sd62;
        fc2_weights[24][30] = 16'sd-20;
        fc2_weights[24][31] = 16'sd18;
        fc2_weights[24][32] = 16'sd-90;
        fc2_weights[24][33] = 16'sd-47;
        fc2_weights[24][34] = 16'sd-37;
        fc2_weights[24][35] = 16'sd-94;
        fc2_weights[24][36] = 16'sd91;
        fc2_weights[24][37] = 16'sd-3;
        fc2_weights[24][38] = 16'sd30;
        fc2_weights[24][39] = 16'sd-27;
        fc2_weights[24][40] = 16'sd-72;
        fc2_weights[24][41] = 16'sd6;
        fc2_weights[24][42] = 16'sd20;
        fc2_weights[24][43] = 16'sd-18;
        fc2_weights[24][44] = 16'sd-12;
        fc2_weights[24][45] = 16'sd16;
        fc2_weights[24][46] = 16'sd14;
        fc2_weights[24][47] = 16'sd-19;
        fc2_weights[24][48] = 16'sd66;
        fc2_weights[24][49] = 16'sd39;
        fc2_weights[24][50] = 16'sd-13;
        fc2_weights[24][51] = 16'sd16;
        fc2_weights[24][52] = 16'sd31;
        fc2_weights[24][53] = 16'sd66;
        fc2_weights[24][54] = 16'sd112;
        fc2_weights[24][55] = 16'sd51;
        fc2_weights[24][56] = 16'sd-22;
        fc2_weights[24][57] = 16'sd-88;
        fc2_weights[24][58] = 16'sd5;
        fc2_weights[24][59] = 16'sd22;
        fc2_weights[24][60] = 16'sd80;
        fc2_weights[24][61] = 16'sd31;
        fc2_weights[24][62] = 16'sd-10;
        fc2_weights[24][63] = 16'sd5;
        fc2_weights[24][64] = 16'sd6;
        fc2_weights[24][65] = 16'sd-28;
        fc2_weights[24][66] = 16'sd-29;
        fc2_weights[24][67] = 16'sd45;
        fc2_weights[24][68] = 16'sd-41;
        fc2_weights[24][69] = 16'sd-17;
        fc2_weights[24][70] = 16'sd67;
        fc2_weights[24][71] = 16'sd-49;
        fc2_weights[24][72] = 16'sd4;
        fc2_weights[24][73] = 16'sd-30;
        fc2_weights[24][74] = 16'sd-13;
        fc2_weights[24][75] = 16'sd14;
        fc2_weights[24][76] = 16'sd-93;
        fc2_weights[24][77] = 16'sd0;
        fc2_weights[24][78] = 16'sd16;
        fc2_weights[24][79] = 16'sd-58;
        fc2_weights[24][80] = 16'sd-48;
        fc2_weights[24][81] = 16'sd82;
        fc2_weights[24][82] = 16'sd5;
        fc2_weights[24][83] = 16'sd-50;
        fc2_weights[24][84] = 16'sd-21;
        fc2_weights[24][85] = 16'sd16;
        fc2_weights[24][86] = 16'sd-25;
        fc2_weights[24][87] = 16'sd-57;
        fc2_weights[24][88] = 16'sd26;
        fc2_weights[24][89] = 16'sd25;
        fc2_weights[24][90] = 16'sd-21;
        fc2_weights[24][91] = 16'sd-18;
        fc2_weights[24][92] = 16'sd34;
        fc2_weights[24][93] = 16'sd13;
        fc2_weights[24][94] = 16'sd-15;
        fc2_weights[24][95] = 16'sd-37;
        fc2_weights[24][96] = 16'sd-79;
        fc2_weights[24][97] = 16'sd24;
        fc2_weights[24][98] = 16'sd14;
        fc2_weights[24][99] = 16'sd28;
        fc2_weights[24][100] = 16'sd31;
        fc2_weights[24][101] = 16'sd-68;
        fc2_weights[24][102] = 16'sd-1;
        fc2_weights[24][103] = 16'sd-52;
        fc2_weights[24][104] = 16'sd-62;
        fc2_weights[24][105] = 16'sd53;
        fc2_weights[24][106] = 16'sd-19;
        fc2_weights[24][107] = 16'sd-29;
        fc2_weights[24][108] = 16'sd27;
        fc2_weights[24][109] = 16'sd40;
        fc2_weights[24][110] = 16'sd-5;
        fc2_weights[24][111] = 16'sd17;
        fc2_weights[24][112] = 16'sd9;
        fc2_weights[24][113] = 16'sd-10;
        fc2_weights[24][114] = 16'sd71;
        fc2_weights[24][115] = 16'sd63;
        fc2_weights[24][116] = 16'sd-45;
        fc2_weights[24][117] = 16'sd-86;
        fc2_weights[24][118] = 16'sd66;
        fc2_weights[24][119] = 16'sd-15;
        fc2_weights[24][120] = 16'sd13;
        fc2_weights[24][121] = 16'sd10;
        fc2_weights[24][122] = 16'sd44;
        fc2_weights[24][123] = 16'sd35;
        fc2_weights[24][124] = 16'sd-37;
        fc2_weights[24][125] = 16'sd-82;
        fc2_weights[24][126] = 16'sd-12;
        fc2_weights[24][127] = 16'sd4;
        fc2_weights[25][0] = 16'sd32;
        fc2_weights[25][1] = 16'sd40;
        fc2_weights[25][2] = 16'sd-84;
        fc2_weights[25][3] = 16'sd55;
        fc2_weights[25][4] = 16'sd-28;
        fc2_weights[25][5] = 16'sd-3;
        fc2_weights[25][6] = 16'sd-4;
        fc2_weights[25][7] = 16'sd2;
        fc2_weights[25][8] = 16'sd1;
        fc2_weights[25][9] = 16'sd35;
        fc2_weights[25][10] = 16'sd-3;
        fc2_weights[25][11] = 16'sd-38;
        fc2_weights[25][12] = 16'sd88;
        fc2_weights[25][13] = 16'sd-20;
        fc2_weights[25][14] = 16'sd1;
        fc2_weights[25][15] = 16'sd-45;
        fc2_weights[25][16] = 16'sd32;
        fc2_weights[25][17] = 16'sd-61;
        fc2_weights[25][18] = 16'sd35;
        fc2_weights[25][19] = 16'sd26;
        fc2_weights[25][20] = 16'sd-65;
        fc2_weights[25][21] = 16'sd-27;
        fc2_weights[25][22] = 16'sd-11;
        fc2_weights[25][23] = 16'sd-17;
        fc2_weights[25][24] = 16'sd-23;
        fc2_weights[25][25] = 16'sd39;
        fc2_weights[25][26] = 16'sd14;
        fc2_weights[25][27] = 16'sd-21;
        fc2_weights[25][28] = 16'sd67;
        fc2_weights[25][29] = 16'sd-13;
        fc2_weights[25][30] = 16'sd-15;
        fc2_weights[25][31] = 16'sd-1;
        fc2_weights[25][32] = 16'sd-17;
        fc2_weights[25][33] = 16'sd8;
        fc2_weights[25][34] = 16'sd1;
        fc2_weights[25][35] = 16'sd-52;
        fc2_weights[25][36] = 16'sd68;
        fc2_weights[25][37] = 16'sd6;
        fc2_weights[25][38] = 16'sd23;
        fc2_weights[25][39] = 16'sd-6;
        fc2_weights[25][40] = 16'sd-44;
        fc2_weights[25][41] = 16'sd3;
        fc2_weights[25][42] = 16'sd-4;
        fc2_weights[25][43] = 16'sd35;
        fc2_weights[25][44] = 16'sd-26;
        fc2_weights[25][45] = 16'sd-76;
        fc2_weights[25][46] = 16'sd-10;
        fc2_weights[25][47] = 16'sd-20;
        fc2_weights[25][48] = 16'sd-55;
        fc2_weights[25][49] = 16'sd-2;
        fc2_weights[25][50] = 16'sd-36;
        fc2_weights[25][51] = 16'sd-42;
        fc2_weights[25][52] = 16'sd-58;
        fc2_weights[25][53] = 16'sd23;
        fc2_weights[25][54] = 16'sd-40;
        fc2_weights[25][55] = 16'sd-11;
        fc2_weights[25][56] = 16'sd-19;
        fc2_weights[25][57] = 16'sd-72;
        fc2_weights[25][58] = 16'sd-21;
        fc2_weights[25][59] = 16'sd42;
        fc2_weights[25][60] = 16'sd-33;
        fc2_weights[25][61] = 16'sd-9;
        fc2_weights[25][62] = 16'sd-88;
        fc2_weights[25][63] = 16'sd-8;
        fc2_weights[25][64] = 16'sd-66;
        fc2_weights[25][65] = 16'sd-34;
        fc2_weights[25][66] = 16'sd-56;
        fc2_weights[25][67] = 16'sd-4;
        fc2_weights[25][68] = 16'sd105;
        fc2_weights[25][69] = 16'sd-37;
        fc2_weights[25][70] = 16'sd-20;
        fc2_weights[25][71] = 16'sd6;
        fc2_weights[25][72] = 16'sd17;
        fc2_weights[25][73] = 16'sd51;
        fc2_weights[25][74] = 16'sd-10;
        fc2_weights[25][75] = 16'sd-2;
        fc2_weights[25][76] = 16'sd-17;
        fc2_weights[25][77] = 16'sd6;
        fc2_weights[25][78] = 16'sd-46;
        fc2_weights[25][79] = 16'sd56;
        fc2_weights[25][80] = 16'sd7;
        fc2_weights[25][81] = 16'sd8;
        fc2_weights[25][82] = 16'sd22;
        fc2_weights[25][83] = 16'sd11;
        fc2_weights[25][84] = 16'sd2;
        fc2_weights[25][85] = 16'sd-50;
        fc2_weights[25][86] = 16'sd-34;
        fc2_weights[25][87] = 16'sd13;
        fc2_weights[25][88] = 16'sd-24;
        fc2_weights[25][89] = 16'sd-41;
        fc2_weights[25][90] = 16'sd-20;
        fc2_weights[25][91] = 16'sd-27;
        fc2_weights[25][92] = 16'sd-26;
        fc2_weights[25][93] = 16'sd22;
        fc2_weights[25][94] = 16'sd20;
        fc2_weights[25][95] = 16'sd-21;
        fc2_weights[25][96] = 16'sd-53;
        fc2_weights[25][97] = 16'sd49;
        fc2_weights[25][98] = 16'sd-18;
        fc2_weights[25][99] = 16'sd21;
        fc2_weights[25][100] = 16'sd-18;
        fc2_weights[25][101] = 16'sd72;
        fc2_weights[25][102] = 16'sd-10;
        fc2_weights[25][103] = 16'sd-97;
        fc2_weights[25][104] = 16'sd-91;
        fc2_weights[25][105] = 16'sd-26;
        fc2_weights[25][106] = 16'sd24;
        fc2_weights[25][107] = 16'sd-44;
        fc2_weights[25][108] = 16'sd19;
        fc2_weights[25][109] = 16'sd7;
        fc2_weights[25][110] = 16'sd-46;
        fc2_weights[25][111] = 16'sd39;
        fc2_weights[25][112] = 16'sd17;
        fc2_weights[25][113] = 16'sd-32;
        fc2_weights[25][114] = 16'sd-20;
        fc2_weights[25][115] = 16'sd29;
        fc2_weights[25][116] = 16'sd15;
        fc2_weights[25][117] = 16'sd-30;
        fc2_weights[25][118] = 16'sd64;
        fc2_weights[25][119] = 16'sd78;
        fc2_weights[25][120] = 16'sd54;
        fc2_weights[25][121] = 16'sd-34;
        fc2_weights[25][122] = 16'sd-90;
        fc2_weights[25][123] = 16'sd-40;
        fc2_weights[25][124] = 16'sd0;
        fc2_weights[25][125] = 16'sd-29;
        fc2_weights[25][126] = 16'sd-24;
        fc2_weights[25][127] = 16'sd-13;
        fc2_weights[26][0] = 16'sd-25;
        fc2_weights[26][1] = 16'sd-8;
        fc2_weights[26][2] = 16'sd15;
        fc2_weights[26][3] = 16'sd5;
        fc2_weights[26][4] = 16'sd6;
        fc2_weights[26][5] = 16'sd32;
        fc2_weights[26][6] = 16'sd-32;
        fc2_weights[26][7] = 16'sd-23;
        fc2_weights[26][8] = 16'sd-52;
        fc2_weights[26][9] = 16'sd35;
        fc2_weights[26][10] = 16'sd-32;
        fc2_weights[26][11] = 16'sd-78;
        fc2_weights[26][12] = 16'sd-3;
        fc2_weights[26][13] = 16'sd39;
        fc2_weights[26][14] = 16'sd8;
        fc2_weights[26][15] = 16'sd-12;
        fc2_weights[26][16] = 16'sd11;
        fc2_weights[26][17] = 16'sd5;
        fc2_weights[26][18] = 16'sd9;
        fc2_weights[26][19] = 16'sd31;
        fc2_weights[26][20] = 16'sd11;
        fc2_weights[26][21] = 16'sd-9;
        fc2_weights[26][22] = 16'sd-14;
        fc2_weights[26][23] = 16'sd-38;
        fc2_weights[26][24] = 16'sd-21;
        fc2_weights[26][25] = 16'sd26;
        fc2_weights[26][26] = 16'sd12;
        fc2_weights[26][27] = 16'sd34;
        fc2_weights[26][28] = 16'sd1;
        fc2_weights[26][29] = 16'sd28;
        fc2_weights[26][30] = 16'sd10;
        fc2_weights[26][31] = 16'sd-10;
        fc2_weights[26][32] = 16'sd-43;
        fc2_weights[26][33] = 16'sd-2;
        fc2_weights[26][34] = 16'sd27;
        fc2_weights[26][35] = 16'sd33;
        fc2_weights[26][36] = 16'sd-16;
        fc2_weights[26][37] = 16'sd-21;
        fc2_weights[26][38] = 16'sd-39;
        fc2_weights[26][39] = 16'sd-40;
        fc2_weights[26][40] = 16'sd34;
        fc2_weights[26][41] = 16'sd-14;
        fc2_weights[26][42] = 16'sd14;
        fc2_weights[26][43] = 16'sd3;
        fc2_weights[26][44] = 16'sd15;
        fc2_weights[26][45] = 16'sd54;
        fc2_weights[26][46] = 16'sd-6;
        fc2_weights[26][47] = 16'sd-30;
        fc2_weights[26][48] = 16'sd61;
        fc2_weights[26][49] = 16'sd17;
        fc2_weights[26][50] = 16'sd29;
        fc2_weights[26][51] = 16'sd1;
        fc2_weights[26][52] = 16'sd22;
        fc2_weights[26][53] = 16'sd-32;
        fc2_weights[26][54] = 16'sd-66;
        fc2_weights[26][55] = 16'sd-17;
        fc2_weights[26][56] = 16'sd24;
        fc2_weights[26][57] = 16'sd-27;
        fc2_weights[26][58] = 16'sd13;
        fc2_weights[26][59] = 16'sd26;
        fc2_weights[26][60] = 16'sd26;
        fc2_weights[26][61] = 16'sd-17;
        fc2_weights[26][62] = 16'sd-13;
        fc2_weights[26][63] = 16'sd5;
        fc2_weights[26][64] = 16'sd-53;
        fc2_weights[26][65] = 16'sd8;
        fc2_weights[26][66] = 16'sd2;
        fc2_weights[26][67] = 16'sd-28;
        fc2_weights[26][68] = 16'sd0;
        fc2_weights[26][69] = 16'sd12;
        fc2_weights[26][70] = 16'sd1;
        fc2_weights[26][71] = 16'sd6;
        fc2_weights[26][72] = 16'sd3;
        fc2_weights[26][73] = 16'sd-63;
        fc2_weights[26][74] = 16'sd-21;
        fc2_weights[26][75] = 16'sd37;
        fc2_weights[26][76] = 16'sd-31;
        fc2_weights[26][77] = 16'sd5;
        fc2_weights[26][78] = 16'sd22;
        fc2_weights[26][79] = 16'sd-18;
        fc2_weights[26][80] = 16'sd-25;
        fc2_weights[26][81] = 16'sd30;
        fc2_weights[26][82] = 16'sd-4;
        fc2_weights[26][83] = 16'sd-24;
        fc2_weights[26][84] = 16'sd4;
        fc2_weights[26][85] = 16'sd18;
        fc2_weights[26][86] = 16'sd-23;
        fc2_weights[26][87] = 16'sd-50;
        fc2_weights[26][88] = 16'sd41;
        fc2_weights[26][89] = 16'sd-68;
        fc2_weights[26][90] = 16'sd19;
        fc2_weights[26][91] = 16'sd-27;
        fc2_weights[26][92] = 16'sd17;
        fc2_weights[26][93] = 16'sd-54;
        fc2_weights[26][94] = 16'sd-28;
        fc2_weights[26][95] = 16'sd-26;
        fc2_weights[26][96] = 16'sd11;
        fc2_weights[26][97] = 16'sd-11;
        fc2_weights[26][98] = 16'sd-19;
        fc2_weights[26][99] = 16'sd-39;
        fc2_weights[26][100] = 16'sd17;
        fc2_weights[26][101] = 16'sd-35;
        fc2_weights[26][102] = 16'sd2;
        fc2_weights[26][103] = 16'sd-10;
        fc2_weights[26][104] = 16'sd33;
        fc2_weights[26][105] = 16'sd11;
        fc2_weights[26][106] = 16'sd23;
        fc2_weights[26][107] = 16'sd19;
        fc2_weights[26][108] = 16'sd-7;
        fc2_weights[26][109] = 16'sd-20;
        fc2_weights[26][110] = 16'sd56;
        fc2_weights[26][111] = 16'sd-18;
        fc2_weights[26][112] = 16'sd-18;
        fc2_weights[26][113] = 16'sd-57;
        fc2_weights[26][114] = 16'sd28;
        fc2_weights[26][115] = 16'sd-26;
        fc2_weights[26][116] = 16'sd-5;
        fc2_weights[26][117] = 16'sd-15;
        fc2_weights[26][118] = 16'sd-16;
        fc2_weights[26][119] = 16'sd-15;
        fc2_weights[26][120] = 16'sd-12;
        fc2_weights[26][121] = 16'sd18;
        fc2_weights[26][122] = 16'sd-4;
        fc2_weights[26][123] = 16'sd66;
        fc2_weights[26][124] = 16'sd-27;
        fc2_weights[26][125] = 16'sd1;
        fc2_weights[26][126] = 16'sd-11;
        fc2_weights[26][127] = 16'sd-70;
        fc2_weights[27][0] = 16'sd39;
        fc2_weights[27][1] = 16'sd2;
        fc2_weights[27][2] = 16'sd-66;
        fc2_weights[27][3] = 16'sd-65;
        fc2_weights[27][4] = 16'sd69;
        fc2_weights[27][5] = 16'sd22;
        fc2_weights[27][6] = 16'sd-5;
        fc2_weights[27][7] = 16'sd-9;
        fc2_weights[27][8] = 16'sd6;
        fc2_weights[27][9] = 16'sd-12;
        fc2_weights[27][10] = 16'sd11;
        fc2_weights[27][11] = 16'sd38;
        fc2_weights[27][12] = 16'sd8;
        fc2_weights[27][13] = 16'sd69;
        fc2_weights[27][14] = 16'sd-33;
        fc2_weights[27][15] = 16'sd18;
        fc2_weights[27][16] = 16'sd-12;
        fc2_weights[27][17] = 16'sd52;
        fc2_weights[27][18] = 16'sd-24;
        fc2_weights[27][19] = 16'sd-18;
        fc2_weights[27][20] = 16'sd2;
        fc2_weights[27][21] = 16'sd-1;
        fc2_weights[27][22] = 16'sd62;
        fc2_weights[27][23] = 16'sd-55;
        fc2_weights[27][24] = 16'sd-10;
        fc2_weights[27][25] = 16'sd-6;
        fc2_weights[27][26] = 16'sd-70;
        fc2_weights[27][27] = 16'sd45;
        fc2_weights[27][28] = 16'sd1;
        fc2_weights[27][29] = 16'sd71;
        fc2_weights[27][30] = 16'sd5;
        fc2_weights[27][31] = 16'sd-8;
        fc2_weights[27][32] = 16'sd-17;
        fc2_weights[27][33] = 16'sd14;
        fc2_weights[27][34] = 16'sd-4;
        fc2_weights[27][35] = 16'sd-26;
        fc2_weights[27][36] = 16'sd-21;
        fc2_weights[27][37] = 16'sd-12;
        fc2_weights[27][38] = 16'sd-34;
        fc2_weights[27][39] = 16'sd-48;
        fc2_weights[27][40] = 16'sd60;
        fc2_weights[27][41] = 16'sd7;
        fc2_weights[27][42] = 16'sd-20;
        fc2_weights[27][43] = 16'sd-11;
        fc2_weights[27][44] = 16'sd-24;
        fc2_weights[27][45] = 16'sd-7;
        fc2_weights[27][46] = 16'sd-67;
        fc2_weights[27][47] = 16'sd-38;
        fc2_weights[27][48] = 16'sd55;
        fc2_weights[27][49] = 16'sd-3;
        fc2_weights[27][50] = 16'sd29;
        fc2_weights[27][51] = 16'sd-12;
        fc2_weights[27][52] = 16'sd15;
        fc2_weights[27][53] = 16'sd-36;
        fc2_weights[27][54] = 16'sd-40;
        fc2_weights[27][55] = 16'sd11;
        fc2_weights[27][56] = 16'sd14;
        fc2_weights[27][57] = 16'sd-57;
        fc2_weights[27][58] = 16'sd11;
        fc2_weights[27][59] = 16'sd-8;
        fc2_weights[27][60] = 16'sd39;
        fc2_weights[27][61] = 16'sd52;
        fc2_weights[27][62] = 16'sd6;
        fc2_weights[27][63] = 16'sd-11;
        fc2_weights[27][64] = 16'sd-30;
        fc2_weights[27][65] = 16'sd-45;
        fc2_weights[27][66] = 16'sd-60;
        fc2_weights[27][67] = 16'sd1;
        fc2_weights[27][68] = 16'sd-9;
        fc2_weights[27][69] = 16'sd-11;
        fc2_weights[27][70] = 16'sd-4;
        fc2_weights[27][71] = 16'sd-43;
        fc2_weights[27][72] = 16'sd-2;
        fc2_weights[27][73] = 16'sd-58;
        fc2_weights[27][74] = 16'sd-26;
        fc2_weights[27][75] = 16'sd12;
        fc2_weights[27][76] = 16'sd-44;
        fc2_weights[27][77] = 16'sd-59;
        fc2_weights[27][78] = 16'sd44;
        fc2_weights[27][79] = 16'sd13;
        fc2_weights[27][80] = 16'sd-25;
        fc2_weights[27][81] = 16'sd-5;
        fc2_weights[27][82] = 16'sd-14;
        fc2_weights[27][83] = 16'sd-17;
        fc2_weights[27][84] = 16'sd-9;
        fc2_weights[27][85] = 16'sd73;
        fc2_weights[27][86] = 16'sd-43;
        fc2_weights[27][87] = 16'sd14;
        fc2_weights[27][88] = 16'sd12;
        fc2_weights[27][89] = 16'sd68;
        fc2_weights[27][90] = 16'sd-38;
        fc2_weights[27][91] = 16'sd-19;
        fc2_weights[27][92] = 16'sd18;
        fc2_weights[27][93] = 16'sd44;
        fc2_weights[27][94] = 16'sd-19;
        fc2_weights[27][95] = 16'sd-24;
        fc2_weights[27][96] = 16'sd-22;
        fc2_weights[27][97] = 16'sd25;
        fc2_weights[27][98] = 16'sd-22;
        fc2_weights[27][99] = 16'sd-6;
        fc2_weights[27][100] = 16'sd-7;
        fc2_weights[27][101] = 16'sd-24;
        fc2_weights[27][102] = 16'sd-53;
        fc2_weights[27][103] = 16'sd14;
        fc2_weights[27][104] = 16'sd1;
        fc2_weights[27][105] = 16'sd39;
        fc2_weights[27][106] = 16'sd-5;
        fc2_weights[27][107] = 16'sd7;
        fc2_weights[27][108] = 16'sd-10;
        fc2_weights[27][109] = 16'sd-72;
        fc2_weights[27][110] = 16'sd41;
        fc2_weights[27][111] = 16'sd-33;
        fc2_weights[27][112] = 16'sd-61;
        fc2_weights[27][113] = 16'sd-27;
        fc2_weights[27][114] = 16'sd11;
        fc2_weights[27][115] = 16'sd6;
        fc2_weights[27][116] = 16'sd2;
        fc2_weights[27][117] = 16'sd27;
        fc2_weights[27][118] = 16'sd0;
        fc2_weights[27][119] = 16'sd-5;
        fc2_weights[27][120] = 16'sd26;
        fc2_weights[27][121] = 16'sd-13;
        fc2_weights[27][122] = 16'sd1;
        fc2_weights[27][123] = 16'sd-24;
        fc2_weights[27][124] = 16'sd-51;
        fc2_weights[27][125] = 16'sd-21;
        fc2_weights[27][126] = 16'sd-23;
        fc2_weights[27][127] = 16'sd48;
        fc2_weights[28][0] = 16'sd-16;
        fc2_weights[28][1] = 16'sd-38;
        fc2_weights[28][2] = 16'sd-39;
        fc2_weights[28][3] = 16'sd-115;
        fc2_weights[28][4] = 16'sd18;
        fc2_weights[28][5] = 16'sd42;
        fc2_weights[28][6] = 16'sd-59;
        fc2_weights[28][7] = 16'sd-31;
        fc2_weights[28][8] = 16'sd1;
        fc2_weights[28][9] = 16'sd-39;
        fc2_weights[28][10] = 16'sd-4;
        fc2_weights[28][11] = 16'sd59;
        fc2_weights[28][12] = 16'sd8;
        fc2_weights[28][13] = 16'sd32;
        fc2_weights[28][14] = 16'sd14;
        fc2_weights[28][15] = 16'sd-36;
        fc2_weights[28][16] = 16'sd0;
        fc2_weights[28][17] = 16'sd-2;
        fc2_weights[28][18] = 16'sd-25;
        fc2_weights[28][19] = 16'sd-50;
        fc2_weights[28][20] = 16'sd8;
        fc2_weights[28][21] = 16'sd6;
        fc2_weights[28][22] = 16'sd23;
        fc2_weights[28][23] = 16'sd-15;
        fc2_weights[28][24] = 16'sd-57;
        fc2_weights[28][25] = 16'sd39;
        fc2_weights[28][26] = 16'sd2;
        fc2_weights[28][27] = 16'sd-23;
        fc2_weights[28][28] = 16'sd-31;
        fc2_weights[28][29] = 16'sd57;
        fc2_weights[28][30] = 16'sd-17;
        fc2_weights[28][31] = 16'sd17;
        fc2_weights[28][32] = 16'sd-66;
        fc2_weights[28][33] = 16'sd-38;
        fc2_weights[28][34] = 16'sd-48;
        fc2_weights[28][35] = 16'sd12;
        fc2_weights[28][36] = 16'sd31;
        fc2_weights[28][37] = 16'sd-49;
        fc2_weights[28][38] = 16'sd57;
        fc2_weights[28][39] = 16'sd36;
        fc2_weights[28][40] = 16'sd-9;
        fc2_weights[28][41] = 16'sd19;
        fc2_weights[28][42] = 16'sd-14;
        fc2_weights[28][43] = 16'sd-30;
        fc2_weights[28][44] = 16'sd-55;
        fc2_weights[28][45] = 16'sd46;
        fc2_weights[28][46] = 16'sd-14;
        fc2_weights[28][47] = 16'sd-59;
        fc2_weights[28][48] = 16'sd75;
        fc2_weights[28][49] = 16'sd56;
        fc2_weights[28][50] = 16'sd54;
        fc2_weights[28][51] = 16'sd39;
        fc2_weights[28][52] = 16'sd-29;
        fc2_weights[28][53] = 16'sd25;
        fc2_weights[28][54] = 16'sd-46;
        fc2_weights[28][55] = 16'sd44;
        fc2_weights[28][56] = 16'sd18;
        fc2_weights[28][57] = 16'sd-44;
        fc2_weights[28][58] = 16'sd-44;
        fc2_weights[28][59] = 16'sd7;
        fc2_weights[28][60] = 16'sd26;
        fc2_weights[28][61] = 16'sd36;
        fc2_weights[28][62] = 16'sd-14;
        fc2_weights[28][63] = 16'sd-108;
        fc2_weights[28][64] = 16'sd-34;
        fc2_weights[28][65] = 16'sd-47;
        fc2_weights[28][66] = 16'sd-24;
        fc2_weights[28][67] = 16'sd8;
        fc2_weights[28][68] = 16'sd-74;
        fc2_weights[28][69] = 16'sd2;
        fc2_weights[28][70] = 16'sd54;
        fc2_weights[28][71] = 16'sd-26;
        fc2_weights[28][72] = 16'sd6;
        fc2_weights[28][73] = 16'sd8;
        fc2_weights[28][74] = 16'sd-61;
        fc2_weights[28][75] = 16'sd53;
        fc2_weights[28][76] = 16'sd-13;
        fc2_weights[28][77] = 16'sd52;
        fc2_weights[28][78] = 16'sd-51;
        fc2_weights[28][79] = 16'sd-14;
        fc2_weights[28][80] = 16'sd-2;
        fc2_weights[28][81] = 16'sd30;
        fc2_weights[28][82] = 16'sd56;
        fc2_weights[28][83] = 16'sd-8;
        fc2_weights[28][84] = 16'sd0;
        fc2_weights[28][85] = 16'sd39;
        fc2_weights[28][86] = 16'sd-37;
        fc2_weights[28][87] = 16'sd-72;
        fc2_weights[28][88] = 16'sd41;
        fc2_weights[28][89] = 16'sd45;
        fc2_weights[28][90] = 16'sd-5;
        fc2_weights[28][91] = 16'sd45;
        fc2_weights[28][92] = 16'sd17;
        fc2_weights[28][93] = 16'sd-38;
        fc2_weights[28][94] = 16'sd-58;
        fc2_weights[28][95] = 16'sd-7;
        fc2_weights[28][96] = 16'sd14;
        fc2_weights[28][97] = 16'sd48;
        fc2_weights[28][98] = 16'sd36;
        fc2_weights[28][99] = 16'sd-34;
        fc2_weights[28][100] = 16'sd39;
        fc2_weights[28][101] = 16'sd-28;
        fc2_weights[28][102] = 16'sd-63;
        fc2_weights[28][103] = 16'sd-3;
        fc2_weights[28][104] = 16'sd-20;
        fc2_weights[28][105] = 16'sd12;
        fc2_weights[28][106] = 16'sd-8;
        fc2_weights[28][107] = 16'sd44;
        fc2_weights[28][108] = 16'sd13;
        fc2_weights[28][109] = 16'sd-12;
        fc2_weights[28][110] = 16'sd-7;
        fc2_weights[28][111] = 16'sd17;
        fc2_weights[28][112] = 16'sd0;
        fc2_weights[28][113] = 16'sd4;
        fc2_weights[28][114] = 16'sd60;
        fc2_weights[28][115] = 16'sd44;
        fc2_weights[28][116] = 16'sd-44;
        fc2_weights[28][117] = 16'sd-37;
        fc2_weights[28][118] = 16'sd83;
        fc2_weights[28][119] = 16'sd-25;
        fc2_weights[28][120] = 16'sd5;
        fc2_weights[28][121] = 16'sd55;
        fc2_weights[28][122] = 16'sd122;
        fc2_weights[28][123] = 16'sd-31;
        fc2_weights[28][124] = 16'sd-23;
        fc2_weights[28][125] = 16'sd-17;
        fc2_weights[28][126] = 16'sd-8;
        fc2_weights[28][127] = 16'sd-31;
        fc2_weights[29][0] = 16'sd-27;
        fc2_weights[29][1] = 16'sd-76;
        fc2_weights[29][2] = 16'sd49;
        fc2_weights[29][3] = 16'sd-40;
        fc2_weights[29][4] = 16'sd-7;
        fc2_weights[29][5] = 16'sd-29;
        fc2_weights[29][6] = 16'sd-23;
        fc2_weights[29][7] = 16'sd11;
        fc2_weights[29][8] = 16'sd9;
        fc2_weights[29][9] = 16'sd-6;
        fc2_weights[29][10] = 16'sd-11;
        fc2_weights[29][11] = 16'sd15;
        fc2_weights[29][12] = 16'sd37;
        fc2_weights[29][13] = 16'sd-7;
        fc2_weights[29][14] = 16'sd-4;
        fc2_weights[29][15] = 16'sd16;
        fc2_weights[29][16] = 16'sd-23;
        fc2_weights[29][17] = 16'sd-20;
        fc2_weights[29][18] = 16'sd-1;
        fc2_weights[29][19] = 16'sd-29;
        fc2_weights[29][20] = 16'sd3;
        fc2_weights[29][21] = 16'sd-19;
        fc2_weights[29][22] = 16'sd-26;
        fc2_weights[29][23] = 16'sd112;
        fc2_weights[29][24] = 16'sd11;
        fc2_weights[29][25] = 16'sd10;
        fc2_weights[29][26] = 16'sd18;
        fc2_weights[29][27] = 16'sd-9;
        fc2_weights[29][28] = 16'sd-62;
        fc2_weights[29][29] = 16'sd8;
        fc2_weights[29][30] = 16'sd-6;
        fc2_weights[29][31] = 16'sd-30;
        fc2_weights[29][32] = 16'sd-24;
        fc2_weights[29][33] = 16'sd-30;
        fc2_weights[29][34] = 16'sd21;
        fc2_weights[29][35] = 16'sd13;
        fc2_weights[29][36] = 16'sd-13;
        fc2_weights[29][37] = 16'sd9;
        fc2_weights[29][38] = 16'sd95;
        fc2_weights[29][39] = 16'sd13;
        fc2_weights[29][40] = 16'sd-49;
        fc2_weights[29][41] = 16'sd-12;
        fc2_weights[29][42] = 16'sd31;
        fc2_weights[29][43] = 16'sd1;
        fc2_weights[29][44] = 16'sd9;
        fc2_weights[29][45] = 16'sd40;
        fc2_weights[29][46] = 16'sd45;
        fc2_weights[29][47] = 16'sd-22;
        fc2_weights[29][48] = 16'sd12;
        fc2_weights[29][49] = 16'sd12;
        fc2_weights[29][50] = 16'sd-1;
        fc2_weights[29][51] = 16'sd-27;
        fc2_weights[29][52] = 16'sd-44;
        fc2_weights[29][53] = 16'sd20;
        fc2_weights[29][54] = 16'sd71;
        fc2_weights[29][55] = 16'sd20;
        fc2_weights[29][56] = 16'sd3;
        fc2_weights[29][57] = 16'sd-19;
        fc2_weights[29][58] = 16'sd45;
        fc2_weights[29][59] = 16'sd0;
        fc2_weights[29][60] = 16'sd-8;
        fc2_weights[29][61] = 16'sd-34;
        fc2_weights[29][62] = 16'sd3;
        fc2_weights[29][63] = 16'sd17;
        fc2_weights[29][64] = 16'sd70;
        fc2_weights[29][65] = 16'sd24;
        fc2_weights[29][66] = 16'sd-43;
        fc2_weights[29][67] = 16'sd12;
        fc2_weights[29][68] = 16'sd-42;
        fc2_weights[29][69] = 16'sd18;
        fc2_weights[29][70] = 16'sd7;
        fc2_weights[29][71] = 16'sd20;
        fc2_weights[29][72] = 16'sd26;
        fc2_weights[29][73] = 16'sd3;
        fc2_weights[29][74] = 16'sd5;
        fc2_weights[29][75] = 16'sd27;
        fc2_weights[29][76] = 16'sd4;
        fc2_weights[29][77] = 16'sd64;
        fc2_weights[29][78] = 16'sd-21;
        fc2_weights[29][79] = 16'sd11;
        fc2_weights[29][80] = 16'sd-71;
        fc2_weights[29][81] = 16'sd9;
        fc2_weights[29][82] = 16'sd-7;
        fc2_weights[29][83] = 16'sd28;
        fc2_weights[29][84] = 16'sd7;
        fc2_weights[29][85] = 16'sd-32;
        fc2_weights[29][86] = 16'sd-9;
        fc2_weights[29][87] = 16'sd-62;
        fc2_weights[29][88] = 16'sd9;
        fc2_weights[29][89] = 16'sd-1;
        fc2_weights[29][90] = 16'sd-22;
        fc2_weights[29][91] = 16'sd-4;
        fc2_weights[29][92] = 16'sd13;
        fc2_weights[29][93] = 16'sd-41;
        fc2_weights[29][94] = 16'sd10;
        fc2_weights[29][95] = 16'sd36;
        fc2_weights[29][96] = 16'sd30;
        fc2_weights[29][97] = 16'sd73;
        fc2_weights[29][98] = 16'sd31;
        fc2_weights[29][99] = 16'sd-14;
        fc2_weights[29][100] = 16'sd19;
        fc2_weights[29][101] = 16'sd-44;
        fc2_weights[29][102] = 16'sd53;
        fc2_weights[29][103] = 16'sd10;
        fc2_weights[29][104] = 16'sd36;
        fc2_weights[29][105] = 16'sd-15;
        fc2_weights[29][106] = 16'sd48;
        fc2_weights[29][107] = 16'sd61;
        fc2_weights[29][108] = 16'sd-54;
        fc2_weights[29][109] = 16'sd-19;
        fc2_weights[29][110] = 16'sd5;
        fc2_weights[29][111] = 16'sd47;
        fc2_weights[29][112] = 16'sd-15;
        fc2_weights[29][113] = 16'sd-17;
        fc2_weights[29][114] = 16'sd55;
        fc2_weights[29][115] = 16'sd-10;
        fc2_weights[29][116] = 16'sd44;
        fc2_weights[29][117] = 16'sd-22;
        fc2_weights[29][118] = 16'sd-5;
        fc2_weights[29][119] = 16'sd-4;
        fc2_weights[29][120] = 16'sd-6;
        fc2_weights[29][121] = 16'sd17;
        fc2_weights[29][122] = 16'sd-12;
        fc2_weights[29][123] = 16'sd28;
        fc2_weights[29][124] = 16'sd38;
        fc2_weights[29][125] = 16'sd5;
        fc2_weights[29][126] = 16'sd18;
        fc2_weights[29][127] = 16'sd-47;
        fc2_weights[30][0] = 16'sd37;
        fc2_weights[30][1] = 16'sd115;
        fc2_weights[30][2] = 16'sd-26;
        fc2_weights[30][3] = 16'sd58;
        fc2_weights[30][4] = 16'sd68;
        fc2_weights[30][5] = 16'sd8;
        fc2_weights[30][6] = 16'sd58;
        fc2_weights[30][7] = 16'sd-5;
        fc2_weights[30][8] = 16'sd18;
        fc2_weights[30][9] = 16'sd-4;
        fc2_weights[30][10] = 16'sd-53;
        fc2_weights[30][11] = 16'sd38;
        fc2_weights[30][12] = 16'sd118;
        fc2_weights[30][13] = 16'sd-7;
        fc2_weights[30][14] = 16'sd-77;
        fc2_weights[30][15] = 16'sd-18;
        fc2_weights[30][16] = 16'sd-70;
        fc2_weights[30][17] = 16'sd42;
        fc2_weights[30][18] = 16'sd-24;
        fc2_weights[30][19] = 16'sd-15;
        fc2_weights[30][20] = 16'sd-8;
        fc2_weights[30][21] = 16'sd2;
        fc2_weights[30][22] = 16'sd5;
        fc2_weights[30][23] = 16'sd-18;
        fc2_weights[30][24] = 16'sd-14;
        fc2_weights[30][25] = 16'sd-37;
        fc2_weights[30][26] = 16'sd0;
        fc2_weights[30][27] = 16'sd-39;
        fc2_weights[30][28] = 16'sd19;
        fc2_weights[30][29] = 16'sd-9;
        fc2_weights[30][30] = 16'sd-7;
        fc2_weights[30][31] = 16'sd15;
        fc2_weights[30][32] = 16'sd27;
        fc2_weights[30][33] = 16'sd42;
        fc2_weights[30][34] = 16'sd-8;
        fc2_weights[30][35] = 16'sd-72;
        fc2_weights[30][36] = 16'sd13;
        fc2_weights[30][37] = 16'sd-26;
        fc2_weights[30][38] = 16'sd25;
        fc2_weights[30][39] = 16'sd45;
        fc2_weights[30][40] = 16'sd-33;
        fc2_weights[30][41] = 16'sd-43;
        fc2_weights[30][42] = 16'sd-43;
        fc2_weights[30][43] = 16'sd32;
        fc2_weights[30][44] = 16'sd-60;
        fc2_weights[30][45] = 16'sd-79;
        fc2_weights[30][46] = 16'sd-52;
        fc2_weights[30][47] = 16'sd42;
        fc2_weights[30][48] = 16'sd-61;
        fc2_weights[30][49] = 16'sd9;
        fc2_weights[30][50] = 16'sd-40;
        fc2_weights[30][51] = 16'sd-98;
        fc2_weights[30][52] = 16'sd-21;
        fc2_weights[30][53] = 16'sd17;
        fc2_weights[30][54] = 16'sd-15;
        fc2_weights[30][55] = 16'sd28;
        fc2_weights[30][56] = 16'sd-2;
        fc2_weights[30][57] = 16'sd-67;
        fc2_weights[30][58] = 16'sd-47;
        fc2_weights[30][59] = 16'sd-55;
        fc2_weights[30][60] = 16'sd-69;
        fc2_weights[30][61] = 16'sd-41;
        fc2_weights[30][62] = 16'sd-92;
        fc2_weights[30][63] = 16'sd-47;
        fc2_weights[30][64] = 16'sd34;
        fc2_weights[30][65] = 16'sd-62;
        fc2_weights[30][66] = 16'sd-88;
        fc2_weights[30][67] = 16'sd-30;
        fc2_weights[30][68] = 16'sd65;
        fc2_weights[30][69] = 16'sd-23;
        fc2_weights[30][70] = 16'sd17;
        fc2_weights[30][71] = 16'sd-43;
        fc2_weights[30][72] = 16'sd68;
        fc2_weights[30][73] = 16'sd10;
        fc2_weights[30][74] = 16'sd-64;
        fc2_weights[30][75] = 16'sd-26;
        fc2_weights[30][76] = 16'sd-45;
        fc2_weights[30][77] = 16'sd-13;
        fc2_weights[30][78] = 16'sd24;
        fc2_weights[30][79] = 16'sd40;
        fc2_weights[30][80] = 16'sd33;
        fc2_weights[30][81] = 16'sd-38;
        fc2_weights[30][82] = 16'sd-51;
        fc2_weights[30][83] = 16'sd-9;
        fc2_weights[30][84] = 16'sd29;
        fc2_weights[30][85] = 16'sd-4;
        fc2_weights[30][86] = 16'sd29;
        fc2_weights[30][87] = 16'sd8;
        fc2_weights[30][88] = 16'sd8;
        fc2_weights[30][89] = 16'sd57;
        fc2_weights[30][90] = 16'sd-84;
        fc2_weights[30][91] = 16'sd-93;
        fc2_weights[30][92] = 16'sd-1;
        fc2_weights[30][93] = 16'sd57;
        fc2_weights[30][94] = 16'sd-23;
        fc2_weights[30][95] = 16'sd9;
        fc2_weights[30][96] = 16'sd-24;
        fc2_weights[30][97] = 16'sd21;
        fc2_weights[30][98] = 16'sd-52;
        fc2_weights[30][99] = 16'sd28;
        fc2_weights[30][100] = 16'sd-82;
        fc2_weights[30][101] = 16'sd48;
        fc2_weights[30][102] = 16'sd-62;
        fc2_weights[30][103] = 16'sd-23;
        fc2_weights[30][104] = 16'sd-48;
        fc2_weights[30][105] = 16'sd-19;
        fc2_weights[30][106] = 16'sd-7;
        fc2_weights[30][107] = 16'sd-12;
        fc2_weights[30][108] = 16'sd-22;
        fc2_weights[30][109] = 16'sd13;
        fc2_weights[30][110] = 16'sd-77;
        fc2_weights[30][111] = 16'sd-57;
        fc2_weights[30][112] = 16'sd44;
        fc2_weights[30][113] = 16'sd3;
        fc2_weights[30][114] = 16'sd-12;
        fc2_weights[30][115] = 16'sd63;
        fc2_weights[30][116] = 16'sd-4;
        fc2_weights[30][117] = 16'sd62;
        fc2_weights[30][118] = 16'sd-5;
        fc2_weights[30][119] = 16'sd45;
        fc2_weights[30][120] = 16'sd22;
        fc2_weights[30][121] = 16'sd-32;
        fc2_weights[30][122] = 16'sd-58;
        fc2_weights[30][123] = 16'sd-72;
        fc2_weights[30][124] = 16'sd-12;
        fc2_weights[30][125] = 16'sd-57;
        fc2_weights[30][126] = 16'sd-60;
        fc2_weights[30][127] = 16'sd4;
        fc2_weights[31][0] = 16'sd-15;
        fc2_weights[31][1] = 16'sd-52;
        fc2_weights[31][2] = 16'sd14;
        fc2_weights[31][3] = 16'sd138;
        fc2_weights[31][4] = 16'sd-11;
        fc2_weights[31][5] = 16'sd-36;
        fc2_weights[31][6] = 16'sd13;
        fc2_weights[31][7] = 16'sd10;
        fc2_weights[31][8] = 16'sd26;
        fc2_weights[31][9] = 16'sd29;
        fc2_weights[31][10] = 16'sd13;
        fc2_weights[31][11] = 16'sd-39;
        fc2_weights[31][12] = 16'sd-7;
        fc2_weights[31][13] = 16'sd1;
        fc2_weights[31][14] = 16'sd25;
        fc2_weights[31][15] = 16'sd62;
        fc2_weights[31][16] = 16'sd-17;
        fc2_weights[31][17] = 16'sd2;
        fc2_weights[31][18] = 16'sd-19;
        fc2_weights[31][19] = 16'sd66;
        fc2_weights[31][20] = 16'sd3;
        fc2_weights[31][21] = 16'sd-37;
        fc2_weights[31][22] = 16'sd-19;
        fc2_weights[31][23] = 16'sd-91;
        fc2_weights[31][24] = 16'sd31;
        fc2_weights[31][25] = 16'sd-56;
        fc2_weights[31][26] = 16'sd69;
        fc2_weights[31][27] = 16'sd-13;
        fc2_weights[31][28] = 16'sd37;
        fc2_weights[31][29] = 16'sd-30;
        fc2_weights[31][30] = 16'sd-11;
        fc2_weights[31][31] = 16'sd6;
        fc2_weights[31][32] = 16'sd-22;
        fc2_weights[31][33] = 16'sd-43;
        fc2_weights[31][34] = 16'sd6;
        fc2_weights[31][35] = 16'sd29;
        fc2_weights[31][36] = 16'sd-46;
        fc2_weights[31][37] = 16'sd-11;
        fc2_weights[31][38] = 16'sd-27;
        fc2_weights[31][39] = 16'sd-48;
        fc2_weights[31][40] = 16'sd-38;
        fc2_weights[31][41] = 16'sd57;
        fc2_weights[31][42] = 16'sd9;
        fc2_weights[31][43] = 16'sd-17;
        fc2_weights[31][44] = 16'sd34;
        fc2_weights[31][45] = 16'sd-41;
        fc2_weights[31][46] = 16'sd13;
        fc2_weights[31][47] = 16'sd7;
        fc2_weights[31][48] = 16'sd-36;
        fc2_weights[31][49] = 16'sd20;
        fc2_weights[31][50] = 16'sd12;
        fc2_weights[31][51] = 16'sd-7;
        fc2_weights[31][52] = 16'sd67;
        fc2_weights[31][53] = 16'sd-12;
        fc2_weights[31][54] = 16'sd-28;
        fc2_weights[31][55] = 16'sd-3;
        fc2_weights[31][56] = 16'sd-15;
        fc2_weights[31][57] = 16'sd-10;
        fc2_weights[31][58] = 16'sd-24;
        fc2_weights[31][59] = 16'sd8;
        fc2_weights[31][60] = 16'sd-22;
        fc2_weights[31][61] = 16'sd5;
        fc2_weights[31][62] = 16'sd27;
        fc2_weights[31][63] = 16'sd23;
        fc2_weights[31][64] = 16'sd-23;
        fc2_weights[31][65] = 16'sd-1;
        fc2_weights[31][66] = 16'sd-26;
        fc2_weights[31][67] = 16'sd20;
        fc2_weights[31][68] = 16'sd43;
        fc2_weights[31][69] = 16'sd-10;
        fc2_weights[31][70] = 16'sd-42;
        fc2_weights[31][71] = 16'sd45;
        fc2_weights[31][72] = 16'sd-25;
        fc2_weights[31][73] = 16'sd35;
        fc2_weights[31][74] = 16'sd-6;
        fc2_weights[31][75] = 16'sd-15;
        fc2_weights[31][76] = 16'sd-3;
        fc2_weights[31][77] = 16'sd-31;
        fc2_weights[31][78] = 16'sd36;
        fc2_weights[31][79] = 16'sd36;
        fc2_weights[31][80] = 16'sd14;
        fc2_weights[31][81] = 16'sd8;
        fc2_weights[31][82] = 16'sd0;
        fc2_weights[31][83] = 16'sd-39;
        fc2_weights[31][84] = 16'sd-15;
        fc2_weights[31][85] = 16'sd-27;
        fc2_weights[31][86] = 16'sd13;
        fc2_weights[31][87] = 16'sd65;
        fc2_weights[31][88] = 16'sd0;
        fc2_weights[31][89] = 16'sd-47;
        fc2_weights[31][90] = 16'sd50;
        fc2_weights[31][91] = 16'sd27;
        fc2_weights[31][92] = 16'sd27;
        fc2_weights[31][93] = 16'sd34;
        fc2_weights[31][94] = 16'sd24;
        fc2_weights[31][95] = 16'sd-1;
        fc2_weights[31][96] = 16'sd3;
        fc2_weights[31][97] = 16'sd-12;
        fc2_weights[31][98] = 16'sd11;
        fc2_weights[31][99] = 16'sd-24;
        fc2_weights[31][100] = 16'sd20;
        fc2_weights[31][101] = 16'sd63;
        fc2_weights[31][102] = 16'sd-33;
        fc2_weights[31][103] = 16'sd-6;
        fc2_weights[31][104] = 16'sd37;
        fc2_weights[31][105] = 16'sd-35;
        fc2_weights[31][106] = 16'sd-9;
        fc2_weights[31][107] = 16'sd32;
        fc2_weights[31][108] = 16'sd3;
        fc2_weights[31][109] = 16'sd37;
        fc2_weights[31][110] = 16'sd-9;
        fc2_weights[31][111] = 16'sd-12;
        fc2_weights[31][112] = 16'sd9;
        fc2_weights[31][113] = 16'sd-12;
        fc2_weights[31][114] = 16'sd5;
        fc2_weights[31][115] = 16'sd-14;
        fc2_weights[31][116] = 16'sd0;
        fc2_weights[31][117] = 16'sd-32;
        fc2_weights[31][118] = 16'sd-57;
        fc2_weights[31][119] = 16'sd-67;
        fc2_weights[31][120] = 16'sd12;
        fc2_weights[31][121] = 16'sd-42;
        fc2_weights[31][122] = 16'sd-3;
        fc2_weights[31][123] = 16'sd-28;
        fc2_weights[31][124] = 16'sd16;
        fc2_weights[31][125] = 16'sd44;
        fc2_weights[31][126] = 16'sd19;
        fc2_weights[31][127] = 16'sd-36;
        fc2_weights[32][0] = 16'sd-12;
        fc2_weights[32][1] = 16'sd32;
        fc2_weights[32][2] = 16'sd-25;
        fc2_weights[32][3] = 16'sd-37;
        fc2_weights[32][4] = 16'sd16;
        fc2_weights[32][5] = 16'sd58;
        fc2_weights[32][6] = 16'sd14;
        fc2_weights[32][7] = 16'sd-2;
        fc2_weights[32][8] = 16'sd129;
        fc2_weights[32][9] = 16'sd17;
        fc2_weights[32][10] = 16'sd-78;
        fc2_weights[32][11] = 16'sd4;
        fc2_weights[32][12] = 16'sd47;
        fc2_weights[32][13] = 16'sd-7;
        fc2_weights[32][14] = 16'sd-78;
        fc2_weights[32][15] = 16'sd-12;
        fc2_weights[32][16] = 16'sd-34;
        fc2_weights[32][17] = 16'sd68;
        fc2_weights[32][18] = 16'sd-37;
        fc2_weights[32][19] = 16'sd-19;
        fc2_weights[32][20] = 16'sd36;
        fc2_weights[32][21] = 16'sd-13;
        fc2_weights[32][22] = 16'sd52;
        fc2_weights[32][23] = 16'sd-6;
        fc2_weights[32][24] = 16'sd-50;
        fc2_weights[32][25] = 16'sd-16;
        fc2_weights[32][26] = 16'sd-67;
        fc2_weights[32][27] = 16'sd-4;
        fc2_weights[32][28] = 16'sd-6;
        fc2_weights[32][29] = 16'sd75;
        fc2_weights[32][30] = 16'sd-12;
        fc2_weights[32][31] = 16'sd-36;
        fc2_weights[32][32] = 16'sd-40;
        fc2_weights[32][33] = 16'sd73;
        fc2_weights[32][34] = 16'sd-4;
        fc2_weights[32][35] = 16'sd-123;
        fc2_weights[32][36] = 16'sd5;
        fc2_weights[32][37] = 16'sd-3;
        fc2_weights[32][38] = 16'sd-14;
        fc2_weights[32][39] = 16'sd42;
        fc2_weights[32][40] = 16'sd2;
        fc2_weights[32][41] = 16'sd75;
        fc2_weights[32][42] = 16'sd15;
        fc2_weights[32][43] = 16'sd20;
        fc2_weights[32][44] = 16'sd-74;
        fc2_weights[32][45] = 16'sd-39;
        fc2_weights[32][46] = 16'sd0;
        fc2_weights[32][47] = 16'sd-10;
        fc2_weights[32][48] = 16'sd-18;
        fc2_weights[32][49] = 16'sd-22;
        fc2_weights[32][50] = 16'sd7;
        fc2_weights[32][51] = 16'sd-25;
        fc2_weights[32][52] = 16'sd-7;
        fc2_weights[32][53] = 16'sd-25;
        fc2_weights[32][54] = 16'sd-4;
        fc2_weights[32][55] = 16'sd6;
        fc2_weights[32][56] = 16'sd3;
        fc2_weights[32][57] = 16'sd-34;
        fc2_weights[32][58] = 16'sd-12;
        fc2_weights[32][59] = 16'sd15;
        fc2_weights[32][60] = 16'sd-1;
        fc2_weights[32][61] = 16'sd41;
        fc2_weights[32][62] = 16'sd-93;
        fc2_weights[32][63] = 16'sd-11;
        fc2_weights[32][64] = 16'sd-41;
        fc2_weights[32][65] = 16'sd-67;
        fc2_weights[32][66] = 16'sd-49;
        fc2_weights[32][67] = 16'sd28;
        fc2_weights[32][68] = 16'sd8;
        fc2_weights[32][69] = 16'sd-15;
        fc2_weights[32][70] = 16'sd22;
        fc2_weights[32][71] = 16'sd-63;
        fc2_weights[32][72] = 16'sd-9;
        fc2_weights[32][73] = 16'sd90;
        fc2_weights[32][74] = 16'sd7;
        fc2_weights[32][75] = 16'sd14;
        fc2_weights[32][76] = 16'sd-28;
        fc2_weights[32][77] = 16'sd30;
        fc2_weights[32][78] = 16'sd-3;
        fc2_weights[32][79] = 16'sd18;
        fc2_weights[32][80] = 16'sd17;
        fc2_weights[32][81] = 16'sd-49;
        fc2_weights[32][82] = 16'sd58;
        fc2_weights[32][83] = 16'sd-69;
        fc2_weights[32][84] = 16'sd35;
        fc2_weights[32][85] = 16'sd62;
        fc2_weights[32][86] = 16'sd-28;
        fc2_weights[32][87] = 16'sd-10;
        fc2_weights[32][88] = 16'sd49;
        fc2_weights[32][89] = 16'sd51;
        fc2_weights[32][90] = 16'sd-1;
        fc2_weights[32][91] = 16'sd-88;
        fc2_weights[32][92] = 16'sd61;
        fc2_weights[32][93] = 16'sd-31;
        fc2_weights[32][94] = 16'sd-6;
        fc2_weights[32][95] = 16'sd-25;
        fc2_weights[32][96] = 16'sd-21;
        fc2_weights[32][97] = 16'sd60;
        fc2_weights[32][98] = 16'sd-41;
        fc2_weights[32][99] = 16'sd-1;
        fc2_weights[32][100] = 16'sd-28;
        fc2_weights[32][101] = 16'sd-44;
        fc2_weights[32][102] = 16'sd-40;
        fc2_weights[32][103] = 16'sd-9;
        fc2_weights[32][104] = 16'sd-52;
        fc2_weights[32][105] = 16'sd-7;
        fc2_weights[32][106] = 16'sd30;
        fc2_weights[32][107] = 16'sd-10;
        fc2_weights[32][108] = 16'sd13;
        fc2_weights[32][109] = 16'sd17;
        fc2_weights[32][110] = 16'sd-4;
        fc2_weights[32][111] = 16'sd37;
        fc2_weights[32][112] = 16'sd14;
        fc2_weights[32][113] = 16'sd74;
        fc2_weights[32][114] = 16'sd59;
        fc2_weights[32][115] = 16'sd61;
        fc2_weights[32][116] = 16'sd-35;
        fc2_weights[32][117] = 16'sd-17;
        fc2_weights[32][118] = 16'sd78;
        fc2_weights[32][119] = 16'sd4;
        fc2_weights[32][120] = 16'sd64;
        fc2_weights[32][121] = 16'sd63;
        fc2_weights[32][122] = 16'sd19;
        fc2_weights[32][123] = 16'sd-53;
        fc2_weights[32][124] = 16'sd41;
        fc2_weights[32][125] = 16'sd-114;
        fc2_weights[32][126] = 16'sd-52;
        fc2_weights[32][127] = 16'sd-24;
        fc2_weights[33][0] = 16'sd-48;
        fc2_weights[33][1] = 16'sd-60;
        fc2_weights[33][2] = 16'sd2;
        fc2_weights[33][3] = 16'sd-33;
        fc2_weights[33][4] = 16'sd13;
        fc2_weights[33][5] = 16'sd34;
        fc2_weights[33][6] = 16'sd-40;
        fc2_weights[33][7] = 16'sd-13;
        fc2_weights[33][8] = 16'sd-56;
        fc2_weights[33][9] = 16'sd14;
        fc2_weights[33][10] = 16'sd2;
        fc2_weights[33][11] = 16'sd-22;
        fc2_weights[33][12] = 16'sd-26;
        fc2_weights[33][13] = 16'sd11;
        fc2_weights[33][14] = 16'sd-15;
        fc2_weights[33][15] = 16'sd15;
        fc2_weights[33][16] = 16'sd11;
        fc2_weights[33][17] = 16'sd34;
        fc2_weights[33][18] = 16'sd6;
        fc2_weights[33][19] = 16'sd21;
        fc2_weights[33][20] = 16'sd-10;
        fc2_weights[33][21] = 16'sd-11;
        fc2_weights[33][22] = 16'sd-12;
        fc2_weights[33][23] = 16'sd-29;
        fc2_weights[33][24] = 16'sd-4;
        fc2_weights[33][25] = 16'sd17;
        fc2_weights[33][26] = 16'sd-41;
        fc2_weights[33][27] = 16'sd41;
        fc2_weights[33][28] = 16'sd-24;
        fc2_weights[33][29] = 16'sd-2;
        fc2_weights[33][30] = 16'sd32;
        fc2_weights[33][31] = 16'sd-28;
        fc2_weights[33][32] = 16'sd-22;
        fc2_weights[33][33] = 16'sd-37;
        fc2_weights[33][34] = 16'sd14;
        fc2_weights[33][35] = 16'sd-6;
        fc2_weights[33][36] = 16'sd-14;
        fc2_weights[33][37] = 16'sd-12;
        fc2_weights[33][38] = 16'sd-13;
        fc2_weights[33][39] = 16'sd-40;
        fc2_weights[33][40] = 16'sd-18;
        fc2_weights[33][41] = 16'sd35;
        fc2_weights[33][42] = 16'sd-21;
        fc2_weights[33][43] = 16'sd-17;
        fc2_weights[33][44] = 16'sd37;
        fc2_weights[33][45] = 16'sd10;
        fc2_weights[33][46] = 16'sd-21;
        fc2_weights[33][47] = 16'sd-17;
        fc2_weights[33][48] = 16'sd60;
        fc2_weights[33][49] = 16'sd19;
        fc2_weights[33][50] = 16'sd41;
        fc2_weights[33][51] = 16'sd17;
        fc2_weights[33][52] = 16'sd9;
        fc2_weights[33][53] = 16'sd-17;
        fc2_weights[33][54] = 16'sd-27;
        fc2_weights[33][55] = 16'sd2;
        fc2_weights[33][56] = 16'sd59;
        fc2_weights[33][57] = 16'sd-28;
        fc2_weights[33][58] = 16'sd8;
        fc2_weights[33][59] = 16'sd23;
        fc2_weights[33][60] = 16'sd36;
        fc2_weights[33][61] = 16'sd-32;
        fc2_weights[33][62] = 16'sd-36;
        fc2_weights[33][63] = 16'sd24;
        fc2_weights[33][64] = 16'sd-57;
        fc2_weights[33][65] = 16'sd-18;
        fc2_weights[33][66] = 16'sd-63;
        fc2_weights[33][67] = 16'sd-32;
        fc2_weights[33][68] = 16'sd-13;
        fc2_weights[33][69] = 16'sd15;
        fc2_weights[33][70] = 16'sd21;
        fc2_weights[33][71] = 16'sd23;
        fc2_weights[33][72] = 16'sd12;
        fc2_weights[33][73] = 16'sd-17;
        fc2_weights[33][74] = 16'sd-37;
        fc2_weights[33][75] = 16'sd8;
        fc2_weights[33][76] = 16'sd12;
        fc2_weights[33][77] = 16'sd49;
        fc2_weights[33][78] = 16'sd6;
        fc2_weights[33][79] = 16'sd-5;
        fc2_weights[33][80] = 16'sd4;
        fc2_weights[33][81] = 16'sd56;
        fc2_weights[33][82] = 16'sd-36;
        fc2_weights[33][83] = 16'sd-22;
        fc2_weights[33][84] = 16'sd-11;
        fc2_weights[33][85] = 16'sd7;
        fc2_weights[33][86] = 16'sd-13;
        fc2_weights[33][87] = 16'sd-9;
        fc2_weights[33][88] = 16'sd61;
        fc2_weights[33][89] = 16'sd-55;
        fc2_weights[33][90] = 16'sd44;
        fc2_weights[33][91] = 16'sd-9;
        fc2_weights[33][92] = 16'sd33;
        fc2_weights[33][93] = 16'sd-38;
        fc2_weights[33][94] = 16'sd-7;
        fc2_weights[33][95] = 16'sd-49;
        fc2_weights[33][96] = 16'sd-2;
        fc2_weights[33][97] = 16'sd-39;
        fc2_weights[33][98] = 16'sd7;
        fc2_weights[33][99] = 16'sd-32;
        fc2_weights[33][100] = 16'sd53;
        fc2_weights[33][101] = 16'sd-44;
        fc2_weights[33][102] = 16'sd54;
        fc2_weights[33][103] = 16'sd120;
        fc2_weights[33][104] = 16'sd11;
        fc2_weights[33][105] = 16'sd-40;
        fc2_weights[33][106] = 16'sd18;
        fc2_weights[33][107] = 16'sd2;
        fc2_weights[33][108] = 16'sd-27;
        fc2_weights[33][109] = 16'sd-37;
        fc2_weights[33][110] = 16'sd11;
        fc2_weights[33][111] = 16'sd-10;
        fc2_weights[33][112] = 16'sd-46;
        fc2_weights[33][113] = 16'sd-6;
        fc2_weights[33][114] = 16'sd6;
        fc2_weights[33][115] = 16'sd-36;
        fc2_weights[33][116] = 16'sd27;
        fc2_weights[33][117] = 16'sd-33;
        fc2_weights[33][118] = 16'sd-53;
        fc2_weights[33][119] = 16'sd-74;
        fc2_weights[33][120] = 16'sd-33;
        fc2_weights[33][121] = 16'sd5;
        fc2_weights[33][122] = 16'sd3;
        fc2_weights[33][123] = 16'sd20;
        fc2_weights[33][124] = 16'sd-17;
        fc2_weights[33][125] = 16'sd-22;
        fc2_weights[33][126] = 16'sd-5;
        fc2_weights[33][127] = 16'sd-13;
        fc2_weights[34][0] = 16'sd-37;
        fc2_weights[34][1] = 16'sd-77;
        fc2_weights[34][2] = 16'sd0;
        fc2_weights[34][3] = 16'sd-68;
        fc2_weights[34][4] = 16'sd16;
        fc2_weights[34][5] = 16'sd8;
        fc2_weights[34][6] = 16'sd-32;
        fc2_weights[34][7] = 16'sd50;
        fc2_weights[34][8] = 16'sd-40;
        fc2_weights[34][9] = 16'sd-33;
        fc2_weights[34][10] = 16'sd58;
        fc2_weights[34][11] = 16'sd-15;
        fc2_weights[34][12] = 16'sd-43;
        fc2_weights[34][13] = 16'sd-21;
        fc2_weights[34][14] = 16'sd-15;
        fc2_weights[34][15] = 16'sd-51;
        fc2_weights[34][16] = 16'sd74;
        fc2_weights[34][17] = 16'sd-83;
        fc2_weights[34][18] = 16'sd-54;
        fc2_weights[34][19] = 16'sd-16;
        fc2_weights[34][20] = 16'sd-87;
        fc2_weights[34][21] = 16'sd50;
        fc2_weights[34][22] = 16'sd24;
        fc2_weights[34][23] = 16'sd38;
        fc2_weights[34][24] = 16'sd57;
        fc2_weights[34][25] = 16'sd27;
        fc2_weights[34][26] = 16'sd20;
        fc2_weights[34][27] = 16'sd-31;
        fc2_weights[34][28] = 16'sd-14;
        fc2_weights[34][29] = 16'sd28;
        fc2_weights[34][30] = 16'sd-38;
        fc2_weights[34][31] = 16'sd-17;
        fc2_weights[34][32] = 16'sd-44;
        fc2_weights[34][33] = 16'sd-57;
        fc2_weights[34][34] = 16'sd3;
        fc2_weights[34][35] = 16'sd7;
        fc2_weights[34][36] = 16'sd-17;
        fc2_weights[34][37] = 16'sd9;
        fc2_weights[34][38] = 16'sd24;
        fc2_weights[34][39] = 16'sd-42;
        fc2_weights[34][40] = 16'sd-17;
        fc2_weights[34][41] = 16'sd12;
        fc2_weights[34][42] = 16'sd13;
        fc2_weights[34][43] = 16'sd-38;
        fc2_weights[34][44] = 16'sd-14;
        fc2_weights[34][45] = 16'sd69;
        fc2_weights[34][46] = 16'sd14;
        fc2_weights[34][47] = 16'sd42;
        fc2_weights[34][48] = 16'sd-76;
        fc2_weights[34][49] = 16'sd-27;
        fc2_weights[34][50] = 16'sd-29;
        fc2_weights[34][51] = 16'sd88;
        fc2_weights[34][52] = 16'sd-58;
        fc2_weights[34][53] = 16'sd21;
        fc2_weights[34][54] = 16'sd49;
        fc2_weights[34][55] = 16'sd11;
        fc2_weights[34][56] = 16'sd8;
        fc2_weights[34][57] = 16'sd-37;
        fc2_weights[34][58] = 16'sd-46;
        fc2_weights[34][59] = 16'sd-6;
        fc2_weights[34][60] = 16'sd81;
        fc2_weights[34][61] = 16'sd46;
        fc2_weights[34][62] = 16'sd-5;
        fc2_weights[34][63] = 16'sd31;
        fc2_weights[34][64] = 16'sd54;
        fc2_weights[34][65] = 16'sd-8;
        fc2_weights[34][66] = 16'sd46;
        fc2_weights[34][67] = 16'sd-17;
        fc2_weights[34][68] = 16'sd-86;
        fc2_weights[34][69] = 16'sd-9;
        fc2_weights[34][70] = 16'sd14;
        fc2_weights[34][71] = 16'sd71;
        fc2_weights[34][72] = 16'sd-36;
        fc2_weights[34][73] = 16'sd-12;
        fc2_weights[34][74] = 16'sd-15;
        fc2_weights[34][75] = 16'sd100;
        fc2_weights[34][76] = 16'sd51;
        fc2_weights[34][77] = 16'sd53;
        fc2_weights[34][78] = 16'sd-75;
        fc2_weights[34][79] = 16'sd18;
        fc2_weights[34][80] = 16'sd3;
        fc2_weights[34][81] = 16'sd-31;
        fc2_weights[34][82] = 16'sd7;
        fc2_weights[34][83] = 16'sd16;
        fc2_weights[34][84] = 16'sd-19;
        fc2_weights[34][85] = 16'sd-12;
        fc2_weights[34][86] = 16'sd8;
        fc2_weights[34][87] = 16'sd-78;
        fc2_weights[34][88] = 16'sd34;
        fc2_weights[34][89] = 16'sd-3;
        fc2_weights[34][90] = 16'sd-18;
        fc2_weights[34][91] = 16'sd9;
        fc2_weights[34][92] = 16'sd64;
        fc2_weights[34][93] = 16'sd5;
        fc2_weights[34][94] = 16'sd-74;
        fc2_weights[34][95] = 16'sd1;
        fc2_weights[34][96] = 16'sd-21;
        fc2_weights[34][97] = 16'sd25;
        fc2_weights[34][98] = 16'sd67;
        fc2_weights[34][99] = 16'sd-61;
        fc2_weights[34][100] = 16'sd21;
        fc2_weights[34][101] = 16'sd-52;
        fc2_weights[34][102] = 16'sd39;
        fc2_weights[34][103] = 16'sd27;
        fc2_weights[34][104] = 16'sd-50;
        fc2_weights[34][105] = 16'sd-16;
        fc2_weights[34][106] = 16'sd14;
        fc2_weights[34][107] = 16'sd-7;
        fc2_weights[34][108] = 16'sd-59;
        fc2_weights[34][109] = 16'sd65;
        fc2_weights[34][110] = 16'sd-21;
        fc2_weights[34][111] = 16'sd38;
        fc2_weights[34][112] = 16'sd-54;
        fc2_weights[34][113] = 16'sd-22;
        fc2_weights[34][114] = 16'sd32;
        fc2_weights[34][115] = 16'sd-41;
        fc2_weights[34][116] = 16'sd35;
        fc2_weights[34][117] = 16'sd-99;
        fc2_weights[34][118] = 16'sd8;
        fc2_weights[34][119] = 16'sd-50;
        fc2_weights[34][120] = 16'sd-20;
        fc2_weights[34][121] = 16'sd44;
        fc2_weights[34][122] = 16'sd37;
        fc2_weights[34][123] = 16'sd-24;
        fc2_weights[34][124] = 16'sd14;
        fc2_weights[34][125] = 16'sd43;
        fc2_weights[34][126] = 16'sd34;
        fc2_weights[34][127] = 16'sd19;
        fc2_weights[35][0] = 16'sd16;
        fc2_weights[35][1] = 16'sd-25;
        fc2_weights[35][2] = 16'sd7;
        fc2_weights[35][3] = 16'sd11;
        fc2_weights[35][4] = 16'sd14;
        fc2_weights[35][5] = 16'sd49;
        fc2_weights[35][6] = 16'sd3;
        fc2_weights[35][7] = 16'sd-15;
        fc2_weights[35][8] = 16'sd-6;
        fc2_weights[35][9] = 16'sd46;
        fc2_weights[35][10] = 16'sd-39;
        fc2_weights[35][11] = 16'sd9;
        fc2_weights[35][12] = 16'sd-8;
        fc2_weights[35][13] = 16'sd79;
        fc2_weights[35][14] = 16'sd26;
        fc2_weights[35][15] = 16'sd3;
        fc2_weights[35][16] = 16'sd19;
        fc2_weights[35][17] = 16'sd74;
        fc2_weights[35][18] = 16'sd30;
        fc2_weights[35][19] = 16'sd-8;
        fc2_weights[35][20] = 16'sd23;
        fc2_weights[35][21] = 16'sd-13;
        fc2_weights[35][22] = 16'sd39;
        fc2_weights[35][23] = 16'sd-19;
        fc2_weights[35][24] = 16'sd-7;
        fc2_weights[35][25] = 16'sd21;
        fc2_weights[35][26] = 16'sd-41;
        fc2_weights[35][27] = 16'sd35;
        fc2_weights[35][28] = 16'sd-5;
        fc2_weights[35][29] = 16'sd11;
        fc2_weights[35][30] = 16'sd56;
        fc2_weights[35][31] = 16'sd-30;
        fc2_weights[35][32] = 16'sd-34;
        fc2_weights[35][33] = 16'sd17;
        fc2_weights[35][34] = 16'sd28;
        fc2_weights[35][35] = 16'sd6;
        fc2_weights[35][36] = 16'sd-5;
        fc2_weights[35][37] = 16'sd-17;
        fc2_weights[35][38] = 16'sd-26;
        fc2_weights[35][39] = 16'sd-44;
        fc2_weights[35][40] = 16'sd25;
        fc2_weights[35][41] = 16'sd-3;
        fc2_weights[35][42] = 16'sd21;
        fc2_weights[35][43] = 16'sd9;
        fc2_weights[35][44] = 16'sd13;
        fc2_weights[35][45] = 16'sd6;
        fc2_weights[35][46] = 16'sd-24;
        fc2_weights[35][47] = 16'sd-6;
        fc2_weights[35][48] = 16'sd61;
        fc2_weights[35][49] = 16'sd-15;
        fc2_weights[35][50] = 16'sd63;
        fc2_weights[35][51] = 16'sd-5;
        fc2_weights[35][52] = 16'sd57;
        fc2_weights[35][53] = 16'sd38;
        fc2_weights[35][54] = 16'sd-42;
        fc2_weights[35][55] = 16'sd19;
        fc2_weights[35][56] = 16'sd37;
        fc2_weights[35][57] = 16'sd-22;
        fc2_weights[35][58] = 16'sd31;
        fc2_weights[35][59] = 16'sd7;
        fc2_weights[35][60] = 16'sd2;
        fc2_weights[35][61] = 16'sd-12;
        fc2_weights[35][62] = 16'sd-14;
        fc2_weights[35][63] = 16'sd1;
        fc2_weights[35][64] = 16'sd-24;
        fc2_weights[35][65] = 16'sd18;
        fc2_weights[35][66] = 16'sd-10;
        fc2_weights[35][67] = 16'sd-2;
        fc2_weights[35][68] = 16'sd-20;
        fc2_weights[35][69] = 16'sd-13;
        fc2_weights[35][70] = 16'sd-1;
        fc2_weights[35][71] = 16'sd-45;
        fc2_weights[35][72] = 16'sd29;
        fc2_weights[35][73] = 16'sd-34;
        fc2_weights[35][74] = 16'sd-7;
        fc2_weights[35][75] = 16'sd33;
        fc2_weights[35][76] = 16'sd-48;
        fc2_weights[35][77] = 16'sd-7;
        fc2_weights[35][78] = 16'sd37;
        fc2_weights[35][79] = 16'sd-33;
        fc2_weights[35][80] = 16'sd-6;
        fc2_weights[35][81] = 16'sd1;
        fc2_weights[35][82] = 16'sd-39;
        fc2_weights[35][83] = 16'sd-14;
        fc2_weights[35][84] = 16'sd-4;
        fc2_weights[35][85] = 16'sd41;
        fc2_weights[35][86] = 16'sd-27;
        fc2_weights[35][87] = 16'sd-31;
        fc2_weights[35][88] = 16'sd20;
        fc2_weights[35][89] = 16'sd-30;
        fc2_weights[35][90] = 16'sd-8;
        fc2_weights[35][91] = 16'sd14;
        fc2_weights[35][92] = 16'sd-14;
        fc2_weights[35][93] = 16'sd-18;
        fc2_weights[35][94] = 16'sd-11;
        fc2_weights[35][95] = 16'sd-20;
        fc2_weights[35][96] = 16'sd-19;
        fc2_weights[35][97] = 16'sd20;
        fc2_weights[35][98] = 16'sd-17;
        fc2_weights[35][99] = 16'sd-16;
        fc2_weights[35][100] = 16'sd-3;
        fc2_weights[35][101] = 16'sd29;
        fc2_weights[35][102] = 16'sd-7;
        fc2_weights[35][103] = 16'sd46;
        fc2_weights[35][104] = 16'sd-20;
        fc2_weights[35][105] = 16'sd36;
        fc2_weights[35][106] = 16'sd7;
        fc2_weights[35][107] = 16'sd12;
        fc2_weights[35][108] = 16'sd5;
        fc2_weights[35][109] = 16'sd-30;
        fc2_weights[35][110] = 16'sd26;
        fc2_weights[35][111] = 16'sd-25;
        fc2_weights[35][112] = 16'sd-13;
        fc2_weights[35][113] = 16'sd-31;
        fc2_weights[35][114] = 16'sd-9;
        fc2_weights[35][115] = 16'sd-26;
        fc2_weights[35][116] = 16'sd1;
        fc2_weights[35][117] = 16'sd15;
        fc2_weights[35][118] = 16'sd-35;
        fc2_weights[35][119] = 16'sd-5;
        fc2_weights[35][120] = 16'sd9;
        fc2_weights[35][121] = 16'sd29;
        fc2_weights[35][122] = 16'sd24;
        fc2_weights[35][123] = 16'sd29;
        fc2_weights[35][124] = 16'sd-30;
        fc2_weights[35][125] = 16'sd-14;
        fc2_weights[35][126] = 16'sd15;
        fc2_weights[35][127] = 16'sd-14;
        fc2_weights[36][0] = 16'sd-69;
        fc2_weights[36][1] = 16'sd92;
        fc2_weights[36][2] = 16'sd-11;
        fc2_weights[36][3] = 16'sd36;
        fc2_weights[36][4] = 16'sd-14;
        fc2_weights[36][5] = 16'sd67;
        fc2_weights[36][6] = 16'sd1;
        fc2_weights[36][7] = 16'sd2;
        fc2_weights[36][8] = 16'sd60;
        fc2_weights[36][9] = 16'sd48;
        fc2_weights[36][10] = 16'sd13;
        fc2_weights[36][11] = 16'sd4;
        fc2_weights[36][12] = 16'sd80;
        fc2_weights[36][13] = 16'sd35;
        fc2_weights[36][14] = 16'sd-48;
        fc2_weights[36][15] = 16'sd-19;
        fc2_weights[36][16] = 16'sd-28;
        fc2_weights[36][17] = 16'sd-59;
        fc2_weights[36][18] = 16'sd44;
        fc2_weights[36][19] = 16'sd11;
        fc2_weights[36][20] = 16'sd-6;
        fc2_weights[36][21] = 16'sd4;
        fc2_weights[36][22] = 16'sd-6;
        fc2_weights[36][23] = 16'sd-29;
        fc2_weights[36][24] = 16'sd1;
        fc2_weights[36][25] = 16'sd-12;
        fc2_weights[36][26] = 16'sd13;
        fc2_weights[36][27] = 16'sd-20;
        fc2_weights[36][28] = 16'sd-14;
        fc2_weights[36][29] = 16'sd-14;
        fc2_weights[36][30] = 16'sd11;
        fc2_weights[36][31] = 16'sd-10;
        fc2_weights[36][32] = 16'sd-5;
        fc2_weights[36][33] = 16'sd29;
        fc2_weights[36][34] = 16'sd-20;
        fc2_weights[36][35] = 16'sd-46;
        fc2_weights[36][36] = 16'sd-4;
        fc2_weights[36][37] = 16'sd55;
        fc2_weights[36][38] = 16'sd-36;
        fc2_weights[36][39] = 16'sd57;
        fc2_weights[36][40] = 16'sd-29;
        fc2_weights[36][41] = 16'sd0;
        fc2_weights[36][42] = 16'sd2;
        fc2_weights[36][43] = 16'sd54;
        fc2_weights[36][44] = 16'sd-3;
        fc2_weights[36][45] = 16'sd-85;
        fc2_weights[36][46] = 16'sd-12;
        fc2_weights[36][47] = 16'sd15;
        fc2_weights[36][48] = 16'sd-22;
        fc2_weights[36][49] = 16'sd-8;
        fc2_weights[36][50] = 16'sd-7;
        fc2_weights[36][51] = 16'sd-58;
        fc2_weights[36][52] = 16'sd-29;
        fc2_weights[36][53] = 16'sd17;
        fc2_weights[36][54] = 16'sd-15;
        fc2_weights[36][55] = 16'sd-28;
        fc2_weights[36][56] = 16'sd22;
        fc2_weights[36][57] = 16'sd-27;
        fc2_weights[36][58] = 16'sd1;
        fc2_weights[36][59] = 16'sd22;
        fc2_weights[36][60] = 16'sd0;
        fc2_weights[36][61] = 16'sd13;
        fc2_weights[36][62] = 16'sd-63;
        fc2_weights[36][63] = 16'sd-8;
        fc2_weights[36][64] = 16'sd-40;
        fc2_weights[36][65] = 16'sd-74;
        fc2_weights[36][66] = 16'sd-6;
        fc2_weights[36][67] = 16'sd-20;
        fc2_weights[36][68] = 16'sd40;
        fc2_weights[36][69] = 16'sd6;
        fc2_weights[36][70] = 16'sd-38;
        fc2_weights[36][71] = 16'sd-9;
        fc2_weights[36][72] = 16'sd62;
        fc2_weights[36][73] = 16'sd18;
        fc2_weights[36][74] = 16'sd0;
        fc2_weights[36][75] = 16'sd-10;
        fc2_weights[36][76] = 16'sd48;
        fc2_weights[36][77] = 16'sd-20;
        fc2_weights[36][78] = 16'sd-43;
        fc2_weights[36][79] = 16'sd27;
        fc2_weights[36][80] = 16'sd24;
        fc2_weights[36][81] = 16'sd-23;
        fc2_weights[36][82] = 16'sd-4;
        fc2_weights[36][83] = 16'sd-19;
        fc2_weights[36][84] = 16'sd4;
        fc2_weights[36][85] = 16'sd0;
        fc2_weights[36][86] = 16'sd-17;
        fc2_weights[36][87] = 16'sd46;
        fc2_weights[36][88] = 16'sd-19;
        fc2_weights[36][89] = 16'sd-15;
        fc2_weights[36][90] = 16'sd-18;
        fc2_weights[36][91] = 16'sd-19;
        fc2_weights[36][92] = 16'sd1;
        fc2_weights[36][93] = 16'sd-16;
        fc2_weights[36][94] = 16'sd41;
        fc2_weights[36][95] = 16'sd-13;
        fc2_weights[36][96] = 16'sd-37;
        fc2_weights[36][97] = 16'sd2;
        fc2_weights[36][98] = 16'sd-18;
        fc2_weights[36][99] = 16'sd-22;
        fc2_weights[36][100] = 16'sd-46;
        fc2_weights[36][101] = 16'sd31;
        fc2_weights[36][102] = 16'sd-24;
        fc2_weights[36][103] = 16'sd-47;
        fc2_weights[36][104] = 16'sd-31;
        fc2_weights[36][105] = 16'sd13;
        fc2_weights[36][106] = 16'sd11;
        fc2_weights[36][107] = 16'sd-25;
        fc2_weights[36][108] = 16'sd19;
        fc2_weights[36][109] = 16'sd14;
        fc2_weights[36][110] = 16'sd-47;
        fc2_weights[36][111] = 16'sd-28;
        fc2_weights[36][112] = 16'sd60;
        fc2_weights[36][113] = 16'sd63;
        fc2_weights[36][114] = 16'sd-6;
        fc2_weights[36][115] = 16'sd18;
        fc2_weights[36][116] = 16'sd-25;
        fc2_weights[36][117] = 16'sd-34;
        fc2_weights[36][118] = 16'sd19;
        fc2_weights[36][119] = 16'sd53;
        fc2_weights[36][120] = 16'sd67;
        fc2_weights[36][121] = 16'sd-21;
        fc2_weights[36][122] = 16'sd-33;
        fc2_weights[36][123] = 16'sd-7;
        fc2_weights[36][124] = 16'sd-21;
        fc2_weights[36][125] = 16'sd-14;
        fc2_weights[36][126] = 16'sd-38;
        fc2_weights[36][127] = 16'sd-68;
        fc2_weights[37][0] = 16'sd-13;
        fc2_weights[37][1] = 16'sd-22;
        fc2_weights[37][2] = 16'sd14;
        fc2_weights[37][3] = 16'sd-7;
        fc2_weights[37][4] = 16'sd-45;
        fc2_weights[37][5] = 16'sd-11;
        fc2_weights[37][6] = 16'sd-27;
        fc2_weights[37][7] = 16'sd11;
        fc2_weights[37][8] = 16'sd-72;
        fc2_weights[37][9] = 16'sd-21;
        fc2_weights[37][10] = 16'sd-39;
        fc2_weights[37][11] = 16'sd-48;
        fc2_weights[37][12] = 16'sd-47;
        fc2_weights[37][13] = 16'sd-20;
        fc2_weights[37][14] = 16'sd29;
        fc2_weights[37][15] = 16'sd21;
        fc2_weights[37][16] = 16'sd1;
        fc2_weights[37][17] = 16'sd-34;
        fc2_weights[37][18] = 16'sd-5;
        fc2_weights[37][19] = 16'sd-31;
        fc2_weights[37][20] = 16'sd-23;
        fc2_weights[37][21] = 16'sd-8;
        fc2_weights[37][22] = 16'sd8;
        fc2_weights[37][23] = 16'sd-5;
        fc2_weights[37][24] = 16'sd19;
        fc2_weights[37][25] = 16'sd-10;
        fc2_weights[37][26] = 16'sd36;
        fc2_weights[37][27] = 16'sd-8;
        fc2_weights[37][28] = 16'sd-31;
        fc2_weights[37][29] = 16'sd-30;
        fc2_weights[37][30] = 16'sd-32;
        fc2_weights[37][31] = 16'sd-9;
        fc2_weights[37][32] = 16'sd-41;
        fc2_weights[37][33] = 16'sd-58;
        fc2_weights[37][34] = 16'sd52;
        fc2_weights[37][35] = 16'sd46;
        fc2_weights[37][36] = 16'sd-18;
        fc2_weights[37][37] = 16'sd-18;
        fc2_weights[37][38] = 16'sd-6;
        fc2_weights[37][39] = 16'sd-35;
        fc2_weights[37][40] = 16'sd-25;
        fc2_weights[37][41] = 16'sd-27;
        fc2_weights[37][42] = 16'sd-12;
        fc2_weights[37][43] = 16'sd-1;
        fc2_weights[37][44] = 16'sd12;
        fc2_weights[37][45] = 16'sd41;
        fc2_weights[37][46] = 16'sd71;
        fc2_weights[37][47] = 16'sd-37;
        fc2_weights[37][48] = 16'sd-31;
        fc2_weights[37][49] = 16'sd19;
        fc2_weights[37][50] = 16'sd-19;
        fc2_weights[37][51] = 16'sd64;
        fc2_weights[37][52] = 16'sd26;
        fc2_weights[37][53] = 16'sd-69;
        fc2_weights[37][54] = 16'sd-10;
        fc2_weights[37][55] = 16'sd-40;
        fc2_weights[37][56] = 16'sd6;
        fc2_weights[37][57] = 16'sd-13;
        fc2_weights[37][58] = 16'sd-8;
        fc2_weights[37][59] = 16'sd-7;
        fc2_weights[37][60] = 16'sd57;
        fc2_weights[37][61] = 16'sd-17;
        fc2_weights[37][62] = 16'sd-4;
        fc2_weights[37][63] = 16'sd5;
        fc2_weights[37][64] = 16'sd26;
        fc2_weights[37][65] = 16'sd33;
        fc2_weights[37][66] = 16'sd29;
        fc2_weights[37][67] = 16'sd-4;
        fc2_weights[37][68] = 16'sd5;
        fc2_weights[37][69] = 16'sd63;
        fc2_weights[37][70] = 16'sd26;
        fc2_weights[37][71] = 16'sd32;
        fc2_weights[37][72] = 16'sd-26;
        fc2_weights[37][73] = 16'sd-22;
        fc2_weights[37][74] = 16'sd8;
        fc2_weights[37][75] = 16'sd-13;
        fc2_weights[37][76] = 16'sd21;
        fc2_weights[37][77] = 16'sd68;
        fc2_weights[37][78] = 16'sd-22;
        fc2_weights[37][79] = 16'sd32;
        fc2_weights[37][80] = 16'sd10;
        fc2_weights[37][81] = 16'sd18;
        fc2_weights[37][82] = 16'sd0;
        fc2_weights[37][83] = 16'sd-2;
        fc2_weights[37][84] = 16'sd-4;
        fc2_weights[37][85] = 16'sd-23;
        fc2_weights[37][86] = 16'sd-25;
        fc2_weights[37][87] = 16'sd-31;
        fc2_weights[37][88] = 16'sd42;
        fc2_weights[37][89] = 16'sd-13;
        fc2_weights[37][90] = 16'sd47;
        fc2_weights[37][91] = 16'sd-32;
        fc2_weights[37][92] = 16'sd41;
        fc2_weights[37][93] = 16'sd-44;
        fc2_weights[37][94] = 16'sd26;
        fc2_weights[37][95] = 16'sd-13;
        fc2_weights[37][96] = 16'sd28;
        fc2_weights[37][97] = 16'sd-48;
        fc2_weights[37][98] = 16'sd-20;
        fc2_weights[37][99] = 16'sd-47;
        fc2_weights[37][100] = 16'sd85;
        fc2_weights[37][101] = 16'sd-75;
        fc2_weights[37][102] = 16'sd40;
        fc2_weights[37][103] = 16'sd-50;
        fc2_weights[37][104] = 16'sd92;
        fc2_weights[37][105] = 16'sd-36;
        fc2_weights[37][106] = 16'sd-15;
        fc2_weights[37][107] = 16'sd9;
        fc2_weights[37][108] = 16'sd-12;
        fc2_weights[37][109] = 16'sd6;
        fc2_weights[37][110] = 16'sd42;
        fc2_weights[37][111] = 16'sd40;
        fc2_weights[37][112] = 16'sd-51;
        fc2_weights[37][113] = 16'sd-54;
        fc2_weights[37][114] = 16'sd10;
        fc2_weights[37][115] = 16'sd-34;
        fc2_weights[37][116] = 16'sd13;
        fc2_weights[37][117] = 16'sd-25;
        fc2_weights[37][118] = 16'sd-37;
        fc2_weights[37][119] = 16'sd-32;
        fc2_weights[37][120] = 16'sd-39;
        fc2_weights[37][121] = 16'sd-53;
        fc2_weights[37][122] = 16'sd46;
        fc2_weights[37][123] = 16'sd0;
        fc2_weights[37][124] = 16'sd-38;
        fc2_weights[37][125] = 16'sd40;
        fc2_weights[37][126] = 16'sd-1;
        fc2_weights[37][127] = 16'sd19;
        fc2_weights[38][0] = 16'sd-45;
        fc2_weights[38][1] = 16'sd6;
        fc2_weights[38][2] = 16'sd3;
        fc2_weights[38][3] = 16'sd47;
        fc2_weights[38][4] = 16'sd-71;
        fc2_weights[38][5] = 16'sd-63;
        fc2_weights[38][6] = 16'sd-64;
        fc2_weights[38][7] = 16'sd-34;
        fc2_weights[38][8] = 16'sd-51;
        fc2_weights[38][9] = 16'sd-2;
        fc2_weights[38][10] = 16'sd7;
        fc2_weights[38][11] = 16'sd1;
        fc2_weights[38][12] = 16'sd-18;
        fc2_weights[38][13] = 16'sd-52;
        fc2_weights[38][14] = 16'sd34;
        fc2_weights[38][15] = 16'sd22;
        fc2_weights[38][16] = 16'sd-41;
        fc2_weights[38][17] = 16'sd-29;
        fc2_weights[38][18] = 16'sd-3;
        fc2_weights[38][19] = 16'sd11;
        fc2_weights[38][20] = 16'sd32;
        fc2_weights[38][21] = 16'sd-26;
        fc2_weights[38][22] = 16'sd-8;
        fc2_weights[38][23] = 16'sd-35;
        fc2_weights[38][24] = 16'sd54;
        fc2_weights[38][25] = 16'sd-23;
        fc2_weights[38][26] = 16'sd53;
        fc2_weights[38][27] = 16'sd-16;
        fc2_weights[38][28] = 16'sd11;
        fc2_weights[38][29] = 16'sd-17;
        fc2_weights[38][30] = 16'sd-28;
        fc2_weights[38][31] = 16'sd-24;
        fc2_weights[38][32] = 16'sd54;
        fc2_weights[38][33] = 16'sd-2;
        fc2_weights[38][34] = 16'sd40;
        fc2_weights[38][35] = 16'sd-20;
        fc2_weights[38][36] = 16'sd-38;
        fc2_weights[38][37] = 16'sd-8;
        fc2_weights[38][38] = 16'sd-33;
        fc2_weights[38][39] = 16'sd0;
        fc2_weights[38][40] = 16'sd-20;
        fc2_weights[38][41] = 16'sd-27;
        fc2_weights[38][42] = 16'sd-21;
        fc2_weights[38][43] = 16'sd-14;
        fc2_weights[38][44] = 16'sd52;
        fc2_weights[38][45] = 16'sd47;
        fc2_weights[38][46] = 16'sd2;
        fc2_weights[38][47] = 16'sd15;
        fc2_weights[38][48] = 16'sd-17;
        fc2_weights[38][49] = 16'sd-17;
        fc2_weights[38][50] = 16'sd-27;
        fc2_weights[38][51] = 16'sd-47;
        fc2_weights[38][52] = 16'sd10;
        fc2_weights[38][53] = 16'sd-25;
        fc2_weights[38][54] = 16'sd-67;
        fc2_weights[38][55] = 16'sd-22;
        fc2_weights[38][56] = 16'sd18;
        fc2_weights[38][57] = 16'sd19;
        fc2_weights[38][58] = 16'sd23;
        fc2_weights[38][59] = 16'sd32;
        fc2_weights[38][60] = 16'sd-8;
        fc2_weights[38][61] = 16'sd6;
        fc2_weights[38][62] = 16'sd-9;
        fc2_weights[38][63] = 16'sd37;
        fc2_weights[38][64] = 16'sd5;
        fc2_weights[38][65] = 16'sd9;
        fc2_weights[38][66] = 16'sd30;
        fc2_weights[38][67] = 16'sd-27;
        fc2_weights[38][68] = 16'sd42;
        fc2_weights[38][69] = 16'sd57;
        fc2_weights[38][70] = 16'sd-39;
        fc2_weights[38][71] = 16'sd42;
        fc2_weights[38][72] = 16'sd-40;
        fc2_weights[38][73] = 16'sd-58;
        fc2_weights[38][74] = 16'sd44;
        fc2_weights[38][75] = 16'sd-29;
        fc2_weights[38][76] = 16'sd-22;
        fc2_weights[38][77] = 16'sd-8;
        fc2_weights[38][78] = 16'sd-38;
        fc2_weights[38][79] = 16'sd28;
        fc2_weights[38][80] = 16'sd-55;
        fc2_weights[38][81] = 16'sd10;
        fc2_weights[38][82] = 16'sd-31;
        fc2_weights[38][83] = 16'sd-25;
        fc2_weights[38][84] = 16'sd-3;
        fc2_weights[38][85] = 16'sd-34;
        fc2_weights[38][86] = 16'sd4;
        fc2_weights[38][87] = 16'sd-9;
        fc2_weights[38][88] = 16'sd49;
        fc2_weights[38][89] = 16'sd-40;
        fc2_weights[38][90] = 16'sd46;
        fc2_weights[38][91] = 16'sd-6;
        fc2_weights[38][92] = 16'sd-1;
        fc2_weights[38][93] = 16'sd-77;
        fc2_weights[38][94] = 16'sd40;
        fc2_weights[38][95] = 16'sd-5;
        fc2_weights[38][96] = 16'sd72;
        fc2_weights[38][97] = 16'sd-39;
        fc2_weights[38][98] = 16'sd27;
        fc2_weights[38][99] = 16'sd-43;
        fc2_weights[38][100] = 16'sd-12;
        fc2_weights[38][101] = 16'sd8;
        fc2_weights[38][102] = 16'sd-6;
        fc2_weights[38][103] = 16'sd-27;
        fc2_weights[38][104] = 16'sd9;
        fc2_weights[38][105] = 16'sd-49;
        fc2_weights[38][106] = 16'sd-22;
        fc2_weights[38][107] = 16'sd63;
        fc2_weights[38][108] = 16'sd6;
        fc2_weights[38][109] = 16'sd-10;
        fc2_weights[38][110] = 16'sd31;
        fc2_weights[38][111] = 16'sd-4;
        fc2_weights[38][112] = 16'sd-25;
        fc2_weights[38][113] = 16'sd-16;
        fc2_weights[38][114] = 16'sd21;
        fc2_weights[38][115] = 16'sd-3;
        fc2_weights[38][116] = 16'sd2;
        fc2_weights[38][117] = 16'sd17;
        fc2_weights[38][118] = 16'sd-34;
        fc2_weights[38][119] = 16'sd14;
        fc2_weights[38][120] = 16'sd-28;
        fc2_weights[38][121] = 16'sd-38;
        fc2_weights[38][122] = 16'sd29;
        fc2_weights[38][123] = 16'sd101;
        fc2_weights[38][124] = 16'sd-9;
        fc2_weights[38][125] = 16'sd31;
        fc2_weights[38][126] = 16'sd-9;
        fc2_weights[38][127] = 16'sd-9;
        fc2_weights[39][0] = 16'sd51;
        fc2_weights[39][1] = 16'sd-18;
        fc2_weights[39][2] = 16'sd-61;
        fc2_weights[39][3] = 16'sd7;
        fc2_weights[39][4] = 16'sd-5;
        fc2_weights[39][5] = 16'sd43;
        fc2_weights[39][6] = 16'sd17;
        fc2_weights[39][7] = 16'sd4;
        fc2_weights[39][8] = 16'sd-21;
        fc2_weights[39][9] = 16'sd-4;
        fc2_weights[39][10] = 16'sd-52;
        fc2_weights[39][11] = 16'sd16;
        fc2_weights[39][12] = 16'sd32;
        fc2_weights[39][13] = 16'sd-11;
        fc2_weights[39][14] = 16'sd5;
        fc2_weights[39][15] = 16'sd-59;
        fc2_weights[39][16] = 16'sd29;
        fc2_weights[39][17] = 16'sd-29;
        fc2_weights[39][18] = 16'sd21;
        fc2_weights[39][19] = 16'sd-27;
        fc2_weights[39][20] = 16'sd33;
        fc2_weights[39][21] = 16'sd-59;
        fc2_weights[39][22] = 16'sd18;
        fc2_weights[39][23] = 16'sd49;
        fc2_weights[39][24] = 16'sd6;
        fc2_weights[39][25] = 16'sd19;
        fc2_weights[39][26] = 16'sd-62;
        fc2_weights[39][27] = 16'sd6;
        fc2_weights[39][28] = 16'sd10;
        fc2_weights[39][29] = 16'sd83;
        fc2_weights[39][30] = 16'sd12;
        fc2_weights[39][31] = 16'sd35;
        fc2_weights[39][32] = 16'sd-36;
        fc2_weights[39][33] = 16'sd19;
        fc2_weights[39][34] = 16'sd-58;
        fc2_weights[39][35] = 16'sd-27;
        fc2_weights[39][36] = 16'sd24;
        fc2_weights[39][37] = 16'sd9;
        fc2_weights[39][38] = 16'sd83;
        fc2_weights[39][39] = 16'sd77;
        fc2_weights[39][40] = 16'sd-37;
        fc2_weights[39][41] = 16'sd-34;
        fc2_weights[39][42] = 16'sd-6;
        fc2_weights[39][43] = 16'sd30;
        fc2_weights[39][44] = 16'sd-54;
        fc2_weights[39][45] = 16'sd-40;
        fc2_weights[39][46] = 16'sd4;
        fc2_weights[39][47] = 16'sd4;
        fc2_weights[39][48] = 16'sd-5;
        fc2_weights[39][49] = 16'sd6;
        fc2_weights[39][50] = 16'sd-5;
        fc2_weights[39][51] = 16'sd-37;
        fc2_weights[39][52] = 16'sd4;
        fc2_weights[39][53] = 16'sd-3;
        fc2_weights[39][54] = 16'sd-42;
        fc2_weights[39][55] = 16'sd4;
        fc2_weights[39][56] = 16'sd-16;
        fc2_weights[39][57] = 16'sd-52;
        fc2_weights[39][58] = 16'sd-19;
        fc2_weights[39][59] = 16'sd-17;
        fc2_weights[39][60] = 16'sd26;
        fc2_weights[39][61] = 16'sd36;
        fc2_weights[39][62] = 16'sd-45;
        fc2_weights[39][63] = 16'sd-1;
        fc2_weights[39][64] = 16'sd-4;
        fc2_weights[39][65] = 16'sd-52;
        fc2_weights[39][66] = 16'sd-16;
        fc2_weights[39][67] = 16'sd47;
        fc2_weights[39][68] = 16'sd-51;
        fc2_weights[39][69] = 16'sd-71;
        fc2_weights[39][70] = 16'sd71;
        fc2_weights[39][71] = 16'sd0;
        fc2_weights[39][72] = 16'sd75;
        fc2_weights[39][73] = 16'sd-42;
        fc2_weights[39][74] = 16'sd-12;
        fc2_weights[39][75] = 16'sd19;
        fc2_weights[39][76] = 16'sd-62;
        fc2_weights[39][77] = 16'sd29;
        fc2_weights[39][78] = 16'sd-37;
        fc2_weights[39][79] = 16'sd-23;
        fc2_weights[39][80] = 16'sd10;
        fc2_weights[39][81] = 16'sd-31;
        fc2_weights[39][82] = 16'sd2;
        fc2_weights[39][83] = 16'sd-29;
        fc2_weights[39][84] = 16'sd-25;
        fc2_weights[39][85] = 16'sd37;
        fc2_weights[39][86] = 16'sd16;
        fc2_weights[39][87] = 16'sd-40;
        fc2_weights[39][88] = 16'sd12;
        fc2_weights[39][89] = 16'sd61;
        fc2_weights[39][90] = 16'sd-55;
        fc2_weights[39][91] = 16'sd-48;
        fc2_weights[39][92] = 16'sd47;
        fc2_weights[39][93] = 16'sd39;
        fc2_weights[39][94] = 16'sd-57;
        fc2_weights[39][95] = 16'sd-48;
        fc2_weights[39][96] = 16'sd-37;
        fc2_weights[39][97] = 16'sd64;
        fc2_weights[39][98] = 16'sd-10;
        fc2_weights[39][99] = 16'sd37;
        fc2_weights[39][100] = 16'sd28;
        fc2_weights[39][101] = 16'sd-25;
        fc2_weights[39][102] = 16'sd-43;
        fc2_weights[39][103] = 16'sd-33;
        fc2_weights[39][104] = 16'sd-7;
        fc2_weights[39][105] = 16'sd38;
        fc2_weights[39][106] = 16'sd-24;
        fc2_weights[39][107] = 16'sd46;
        fc2_weights[39][108] = 16'sd56;
        fc2_weights[39][109] = 16'sd33;
        fc2_weights[39][110] = 16'sd-14;
        fc2_weights[39][111] = 16'sd-37;
        fc2_weights[39][112] = 16'sd19;
        fc2_weights[39][113] = 16'sd-23;
        fc2_weights[39][114] = 16'sd80;
        fc2_weights[39][115] = 16'sd58;
        fc2_weights[39][116] = 16'sd-40;
        fc2_weights[39][117] = 16'sd-15;
        fc2_weights[39][118] = 16'sd62;
        fc2_weights[39][119] = 16'sd-3;
        fc2_weights[39][120] = 16'sd-6;
        fc2_weights[39][121] = 16'sd38;
        fc2_weights[39][122] = 16'sd-1;
        fc2_weights[39][123] = 16'sd-50;
        fc2_weights[39][124] = 16'sd14;
        fc2_weights[39][125] = 16'sd-55;
        fc2_weights[39][126] = 16'sd-36;
        fc2_weights[39][127] = 16'sd-29;
        fc2_weights[40][0] = 16'sd35;
        fc2_weights[40][1] = 16'sd-32;
        fc2_weights[40][2] = 16'sd41;
        fc2_weights[40][3] = 16'sd-32;
        fc2_weights[40][4] = 16'sd21;
        fc2_weights[40][5] = 16'sd-20;
        fc2_weights[40][6] = 16'sd-11;
        fc2_weights[40][7] = 16'sd23;
        fc2_weights[40][8] = 16'sd-40;
        fc2_weights[40][9] = 16'sd72;
        fc2_weights[40][10] = 16'sd-57;
        fc2_weights[40][11] = 16'sd3;
        fc2_weights[40][12] = 16'sd-6;
        fc2_weights[40][13] = 16'sd11;
        fc2_weights[40][14] = 16'sd24;
        fc2_weights[40][15] = 16'sd-6;
        fc2_weights[40][16] = 16'sd-38;
        fc2_weights[40][17] = 16'sd-18;
        fc2_weights[40][18] = 16'sd116;
        fc2_weights[40][19] = 16'sd-19;
        fc2_weights[40][20] = 16'sd20;
        fc2_weights[40][21] = 16'sd-34;
        fc2_weights[40][22] = 16'sd15;
        fc2_weights[40][23] = 16'sd0;
        fc2_weights[40][24] = 16'sd-27;
        fc2_weights[40][25] = 16'sd9;
        fc2_weights[40][26] = 16'sd33;
        fc2_weights[40][27] = 16'sd50;
        fc2_weights[40][28] = 16'sd-39;
        fc2_weights[40][29] = 16'sd40;
        fc2_weights[40][30] = 16'sd0;
        fc2_weights[40][31] = 16'sd13;
        fc2_weights[40][32] = 16'sd-56;
        fc2_weights[40][33] = 16'sd-30;
        fc2_weights[40][34] = 16'sd-9;
        fc2_weights[40][35] = 16'sd-37;
        fc2_weights[40][36] = 16'sd4;
        fc2_weights[40][37] = 16'sd54;
        fc2_weights[40][38] = 16'sd67;
        fc2_weights[40][39] = 16'sd6;
        fc2_weights[40][40] = 16'sd-43;
        fc2_weights[40][41] = 16'sd31;
        fc2_weights[40][42] = 16'sd51;
        fc2_weights[40][43] = 16'sd31;
        fc2_weights[40][44] = 16'sd-27;
        fc2_weights[40][45] = 16'sd50;
        fc2_weights[40][46] = 16'sd11;
        fc2_weights[40][47] = 16'sd-20;
        fc2_weights[40][48] = 16'sd-14;
        fc2_weights[40][49] = 16'sd9;
        fc2_weights[40][50] = 16'sd35;
        fc2_weights[40][51] = 16'sd-10;
        fc2_weights[40][52] = 16'sd42;
        fc2_weights[40][53] = 16'sd42;
        fc2_weights[40][54] = 16'sd-5;
        fc2_weights[40][55] = 16'sd4;
        fc2_weights[40][56] = 16'sd10;
        fc2_weights[40][57] = 16'sd-63;
        fc2_weights[40][58] = 16'sd38;
        fc2_weights[40][59] = 16'sd-28;
        fc2_weights[40][60] = 16'sd-29;
        fc2_weights[40][61] = 16'sd17;
        fc2_weights[40][62] = 16'sd30;
        fc2_weights[40][63] = 16'sd20;
        fc2_weights[40][64] = 16'sd1;
        fc2_weights[40][65] = 16'sd53;
        fc2_weights[40][66] = 16'sd-25;
        fc2_weights[40][67] = 16'sd72;
        fc2_weights[40][68] = 16'sd0;
        fc2_weights[40][69] = 16'sd-54;
        fc2_weights[40][70] = 16'sd3;
        fc2_weights[40][71] = 16'sd-40;
        fc2_weights[40][72] = 16'sd55;
        fc2_weights[40][73] = 16'sd8;
        fc2_weights[40][74] = 16'sd39;
        fc2_weights[40][75] = 16'sd10;
        fc2_weights[40][76] = 16'sd-68;
        fc2_weights[40][77] = 16'sd12;
        fc2_weights[40][78] = 16'sd9;
        fc2_weights[40][79] = 16'sd1;
        fc2_weights[40][80] = 16'sd-62;
        fc2_weights[40][81] = 16'sd31;
        fc2_weights[40][82] = 16'sd26;
        fc2_weights[40][83] = 16'sd-65;
        fc2_weights[40][84] = 16'sd35;
        fc2_weights[40][85] = 16'sd5;
        fc2_weights[40][86] = 16'sd-27;
        fc2_weights[40][87] = 16'sd-27;
        fc2_weights[40][88] = 16'sd-22;
        fc2_weights[40][89] = 16'sd33;
        fc2_weights[40][90] = 16'sd18;
        fc2_weights[40][91] = 16'sd28;
        fc2_weights[40][92] = 16'sd0;
        fc2_weights[40][93] = 16'sd-71;
        fc2_weights[40][94] = 16'sd-1;
        fc2_weights[40][95] = 16'sd-3;
        fc2_weights[40][96] = 16'sd-32;
        fc2_weights[40][97] = 16'sd78;
        fc2_weights[40][98] = 16'sd-2;
        fc2_weights[40][99] = 16'sd96;
        fc2_weights[40][100] = 16'sd67;
        fc2_weights[40][101] = 16'sd11;
        fc2_weights[40][102] = 16'sd16;
        fc2_weights[40][103] = 16'sd-31;
        fc2_weights[40][104] = 16'sd36;
        fc2_weights[40][105] = 16'sd20;
        fc2_weights[40][106] = 16'sd32;
        fc2_weights[40][107] = 16'sd41;
        fc2_weights[40][108] = 16'sd45;
        fc2_weights[40][109] = 16'sd-30;
        fc2_weights[40][110] = 16'sd17;
        fc2_weights[40][111] = 16'sd1;
        fc2_weights[40][112] = 16'sd16;
        fc2_weights[40][113] = 16'sd3;
        fc2_weights[40][114] = 16'sd33;
        fc2_weights[40][115] = 16'sd-5;
        fc2_weights[40][116] = 16'sd8;
        fc2_weights[40][117] = 16'sd-39;
        fc2_weights[40][118] = 16'sd19;
        fc2_weights[40][119] = 16'sd-38;
        fc2_weights[40][120] = 16'sd-29;
        fc2_weights[40][121] = 16'sd27;
        fc2_weights[40][122] = 16'sd41;
        fc2_weights[40][123] = 16'sd23;
        fc2_weights[40][124] = 16'sd-19;
        fc2_weights[40][125] = 16'sd-9;
        fc2_weights[40][126] = 16'sd-2;
        fc2_weights[40][127] = 16'sd-37;
        fc2_weights[41][0] = 16'sd-27;
        fc2_weights[41][1] = 16'sd-2;
        fc2_weights[41][2] = 16'sd-17;
        fc2_weights[41][3] = 16'sd0;
        fc2_weights[41][4] = 16'sd-7;
        fc2_weights[41][5] = 16'sd14;
        fc2_weights[41][6] = 16'sd28;
        fc2_weights[41][7] = 16'sd10;
        fc2_weights[41][8] = 16'sd15;
        fc2_weights[41][9] = 16'sd-10;
        fc2_weights[41][10] = 16'sd-32;
        fc2_weights[41][11] = 16'sd2;
        fc2_weights[41][12] = 16'sd-44;
        fc2_weights[41][13] = 16'sd30;
        fc2_weights[41][14] = 16'sd61;
        fc2_weights[41][15] = 16'sd-11;
        fc2_weights[41][16] = 16'sd-21;
        fc2_weights[41][17] = 16'sd12;
        fc2_weights[41][18] = 16'sd-21;
        fc2_weights[41][19] = 16'sd67;
        fc2_weights[41][20] = 16'sd39;
        fc2_weights[41][21] = 16'sd-5;
        fc2_weights[41][22] = 16'sd45;
        fc2_weights[41][23] = 16'sd-54;
        fc2_weights[41][24] = 16'sd11;
        fc2_weights[41][25] = 16'sd2;
        fc2_weights[41][26] = 16'sd-22;
        fc2_weights[41][27] = 16'sd-11;
        fc2_weights[41][28] = 16'sd9;
        fc2_weights[41][29] = 16'sd11;
        fc2_weights[41][30] = 16'sd-10;
        fc2_weights[41][31] = 16'sd-20;
        fc2_weights[41][32] = 16'sd-36;
        fc2_weights[41][33] = 16'sd-37;
        fc2_weights[41][34] = 16'sd25;
        fc2_weights[41][35] = 16'sd-14;
        fc2_weights[41][36] = 16'sd-28;
        fc2_weights[41][37] = 16'sd-21;
        fc2_weights[41][38] = 16'sd27;
        fc2_weights[41][39] = 16'sd-11;
        fc2_weights[41][40] = 16'sd-31;
        fc2_weights[41][41] = 16'sd-32;
        fc2_weights[41][42] = 16'sd4;
        fc2_weights[41][43] = 16'sd-23;
        fc2_weights[41][44] = 16'sd-10;
        fc2_weights[41][45] = 16'sd3;
        fc2_weights[41][46] = 16'sd12;
        fc2_weights[41][47] = 16'sd28;
        fc2_weights[41][48] = 16'sd-3;
        fc2_weights[41][49] = 16'sd23;
        fc2_weights[41][50] = 16'sd-21;
        fc2_weights[41][51] = 16'sd-6;
        fc2_weights[41][52] = 16'sd101;
        fc2_weights[41][53] = 16'sd-50;
        fc2_weights[41][54] = 16'sd22;
        fc2_weights[41][55] = 16'sd-34;
        fc2_weights[41][56] = 16'sd0;
        fc2_weights[41][57] = 16'sd-6;
        fc2_weights[41][58] = 16'sd-3;
        fc2_weights[41][59] = 16'sd57;
        fc2_weights[41][60] = 16'sd11;
        fc2_weights[41][61] = 16'sd-41;
        fc2_weights[41][62] = 16'sd71;
        fc2_weights[41][63] = 16'sd-5;
        fc2_weights[41][64] = 16'sd-7;
        fc2_weights[41][65] = 16'sd44;
        fc2_weights[41][66] = 16'sd2;
        fc2_weights[41][67] = 16'sd51;
        fc2_weights[41][68] = 16'sd14;
        fc2_weights[41][69] = 16'sd-5;
        fc2_weights[41][70] = 16'sd-45;
        fc2_weights[41][71] = 16'sd0;
        fc2_weights[41][72] = 16'sd-9;
        fc2_weights[41][73] = 16'sd-19;
        fc2_weights[41][74] = 16'sd-11;
        fc2_weights[41][75] = 16'sd-20;
        fc2_weights[41][76] = 16'sd-51;
        fc2_weights[41][77] = 16'sd-19;
        fc2_weights[41][78] = 16'sd-45;
        fc2_weights[41][79] = 16'sd31;
        fc2_weights[41][80] = 16'sd13;
        fc2_weights[41][81] = 16'sd21;
        fc2_weights[41][82] = 16'sd26;
        fc2_weights[41][83] = 16'sd-73;
        fc2_weights[41][84] = 16'sd22;
        fc2_weights[41][85] = 16'sd9;
        fc2_weights[41][86] = 16'sd-24;
        fc2_weights[41][87] = 16'sd-9;
        fc2_weights[41][88] = 16'sd7;
        fc2_weights[41][89] = 16'sd17;
        fc2_weights[41][90] = 16'sd67;
        fc2_weights[41][91] = 16'sd-31;
        fc2_weights[41][92] = 16'sd43;
        fc2_weights[41][93] = 16'sd36;
        fc2_weights[41][94] = 16'sd-39;
        fc2_weights[41][95] = 16'sd-8;
        fc2_weights[41][96] = 16'sd-46;
        fc2_weights[41][97] = 16'sd6;
        fc2_weights[41][98] = 16'sd-13;
        fc2_weights[41][99] = 16'sd-1;
        fc2_weights[41][100] = 16'sd15;
        fc2_weights[41][101] = 16'sd-8;
        fc2_weights[41][102] = 16'sd-34;
        fc2_weights[41][103] = 16'sd-29;
        fc2_weights[41][104] = 16'sd-16;
        fc2_weights[41][105] = 16'sd-23;
        fc2_weights[41][106] = 16'sd-26;
        fc2_weights[41][107] = 16'sd-21;
        fc2_weights[41][108] = 16'sd-24;
        fc2_weights[41][109] = 16'sd16;
        fc2_weights[41][110] = 16'sd-37;
        fc2_weights[41][111] = 16'sd-15;
        fc2_weights[41][112] = 16'sd-45;
        fc2_weights[41][113] = 16'sd-31;
        fc2_weights[41][114] = 16'sd11;
        fc2_weights[41][115] = 16'sd14;
        fc2_weights[41][116] = 16'sd-11;
        fc2_weights[41][117] = 16'sd29;
        fc2_weights[41][118] = 16'sd25;
        fc2_weights[41][119] = 16'sd-58;
        fc2_weights[41][120] = 16'sd-32;
        fc2_weights[41][121] = 16'sd-32;
        fc2_weights[41][122] = 16'sd-88;
        fc2_weights[41][123] = 16'sd-31;
        fc2_weights[41][124] = 16'sd8;
        fc2_weights[41][125] = 16'sd-14;
        fc2_weights[41][126] = 16'sd36;
        fc2_weights[41][127] = 16'sd75;
        fc2_weights[42][0] = 16'sd5;
        fc2_weights[42][1] = 16'sd-11;
        fc2_weights[42][2] = 16'sd-29;
        fc2_weights[42][3] = 16'sd-2;
        fc2_weights[42][4] = 16'sd36;
        fc2_weights[42][5] = 16'sd2;
        fc2_weights[42][6] = 16'sd30;
        fc2_weights[42][7] = 16'sd-17;
        fc2_weights[42][8] = 16'sd0;
        fc2_weights[42][9] = 16'sd-29;
        fc2_weights[42][10] = 16'sd-21;
        fc2_weights[42][11] = 16'sd11;
        fc2_weights[42][12] = 16'sd27;
        fc2_weights[42][13] = 16'sd33;
        fc2_weights[42][14] = 16'sd-3;
        fc2_weights[42][15] = 16'sd4;
        fc2_weights[42][16] = 16'sd-47;
        fc2_weights[42][17] = 16'sd81;
        fc2_weights[42][18] = 16'sd-7;
        fc2_weights[42][19] = 16'sd18;
        fc2_weights[42][20] = 16'sd56;
        fc2_weights[42][21] = 16'sd-26;
        fc2_weights[42][22] = 16'sd41;
        fc2_weights[42][23] = 16'sd-27;
        fc2_weights[42][24] = 16'sd40;
        fc2_weights[42][25] = 16'sd-26;
        fc2_weights[42][26] = 16'sd-65;
        fc2_weights[42][27] = 16'sd-15;
        fc2_weights[42][28] = 16'sd-8;
        fc2_weights[42][29] = 16'sd15;
        fc2_weights[42][30] = 16'sd34;
        fc2_weights[42][31] = 16'sd8;
        fc2_weights[42][32] = 16'sd20;
        fc2_weights[42][33] = 16'sd29;
        fc2_weights[42][34] = 16'sd-22;
        fc2_weights[42][35] = 16'sd8;
        fc2_weights[42][36] = 16'sd-5;
        fc2_weights[42][37] = 16'sd-29;
        fc2_weights[42][38] = 16'sd-41;
        fc2_weights[42][39] = 16'sd-15;
        fc2_weights[42][40] = 16'sd58;
        fc2_weights[42][41] = 16'sd-71;
        fc2_weights[42][42] = 16'sd45;
        fc2_weights[42][43] = 16'sd16;
        fc2_weights[42][44] = 16'sd-5;
        fc2_weights[42][45] = 16'sd5;
        fc2_weights[42][46] = 16'sd-35;
        fc2_weights[42][47] = 16'sd5;
        fc2_weights[42][48] = 16'sd-9;
        fc2_weights[42][49] = 16'sd-25;
        fc2_weights[42][50] = 16'sd15;
        fc2_weights[42][51] = 16'sd14;
        fc2_weights[42][52] = 16'sd52;
        fc2_weights[42][53] = 16'sd10;
        fc2_weights[42][54] = 16'sd-73;
        fc2_weights[42][55] = 16'sd-5;
        fc2_weights[42][56] = 16'sd-3;
        fc2_weights[42][57] = 16'sd-18;
        fc2_weights[42][58] = 16'sd43;
        fc2_weights[42][59] = 16'sd62;
        fc2_weights[42][60] = 16'sd17;
        fc2_weights[42][61] = 16'sd10;
        fc2_weights[42][62] = 16'sd33;
        fc2_weights[42][63] = 16'sd9;
        fc2_weights[42][64] = 16'sd-42;
        fc2_weights[42][65] = 16'sd-11;
        fc2_weights[42][66] = 16'sd-61;
        fc2_weights[42][67] = 16'sd3;
        fc2_weights[42][68] = 16'sd-55;
        fc2_weights[42][69] = 16'sd45;
        fc2_weights[42][70] = 16'sd-63;
        fc2_weights[42][71] = 16'sd-43;
        fc2_weights[42][72] = 16'sd3;
        fc2_weights[42][73] = 16'sd-45;
        fc2_weights[42][74] = 16'sd-16;
        fc2_weights[42][75] = 16'sd-33;
        fc2_weights[42][76] = 16'sd-55;
        fc2_weights[42][77] = 16'sd-72;
        fc2_weights[42][78] = 16'sd54;
        fc2_weights[42][79] = 16'sd-38;
        fc2_weights[42][80] = 16'sd-42;
        fc2_weights[42][81] = 16'sd-19;
        fc2_weights[42][82] = 16'sd11;
        fc2_weights[42][83] = 16'sd-44;
        fc2_weights[42][84] = 16'sd15;
        fc2_weights[42][85] = 16'sd-2;
        fc2_weights[42][86] = 16'sd-49;
        fc2_weights[42][87] = 16'sd30;
        fc2_weights[42][88] = 16'sd5;
        fc2_weights[42][89] = 16'sd-29;
        fc2_weights[42][90] = 16'sd8;
        fc2_weights[42][91] = 16'sd-38;
        fc2_weights[42][92] = 16'sd-31;
        fc2_weights[42][93] = 16'sd23;
        fc2_weights[42][94] = 16'sd-39;
        fc2_weights[42][95] = 16'sd-24;
        fc2_weights[42][96] = 16'sd26;
        fc2_weights[42][97] = 16'sd9;
        fc2_weights[42][98] = 16'sd-45;
        fc2_weights[42][99] = 16'sd-13;
        fc2_weights[42][100] = 16'sd13;
        fc2_weights[42][101] = 16'sd8;
        fc2_weights[42][102] = 16'sd-12;
        fc2_weights[42][103] = 16'sd67;
        fc2_weights[42][104] = 16'sd-18;
        fc2_weights[42][105] = 16'sd8;
        fc2_weights[42][106] = 16'sd-10;
        fc2_weights[42][107] = 16'sd-46;
        fc2_weights[42][108] = 16'sd-32;
        fc2_weights[42][109] = 16'sd-68;
        fc2_weights[42][110] = 16'sd4;
        fc2_weights[42][111] = 16'sd-39;
        fc2_weights[42][112] = 16'sd-68;
        fc2_weights[42][113] = 16'sd-13;
        fc2_weights[42][114] = 16'sd-7;
        fc2_weights[42][115] = 16'sd-29;
        fc2_weights[42][116] = 16'sd0;
        fc2_weights[42][117] = 16'sd65;
        fc2_weights[42][118] = 16'sd-72;
        fc2_weights[42][119] = 16'sd19;
        fc2_weights[42][120] = 16'sd14;
        fc2_weights[42][121] = 16'sd-61;
        fc2_weights[42][122] = 16'sd-22;
        fc2_weights[42][123] = 16'sd7;
        fc2_weights[42][124] = 16'sd13;
        fc2_weights[42][125] = 16'sd8;
        fc2_weights[42][126] = 16'sd43;
        fc2_weights[42][127] = 16'sd55;
        fc2_weights[43][0] = 16'sd-21;
        fc2_weights[43][1] = 16'sd13;
        fc2_weights[43][2] = 16'sd-30;
        fc2_weights[43][3] = 16'sd-51;
        fc2_weights[43][4] = 16'sd60;
        fc2_weights[43][5] = 16'sd42;
        fc2_weights[43][6] = 16'sd-12;
        fc2_weights[43][7] = 16'sd23;
        fc2_weights[43][8] = 16'sd-6;
        fc2_weights[43][9] = 16'sd-22;
        fc2_weights[43][10] = 16'sd44;
        fc2_weights[43][11] = 16'sd6;
        fc2_weights[43][12] = 16'sd22;
        fc2_weights[43][13] = 16'sd15;
        fc2_weights[43][14] = 16'sd-31;
        fc2_weights[43][15] = 16'sd-30;
        fc2_weights[43][16] = 16'sd-7;
        fc2_weights[43][17] = 16'sd-29;
        fc2_weights[43][18] = 16'sd-74;
        fc2_weights[43][19] = 16'sd-59;
        fc2_weights[43][20] = 16'sd21;
        fc2_weights[43][21] = 16'sd6;
        fc2_weights[43][22] = 16'sd56;
        fc2_weights[43][23] = 16'sd22;
        fc2_weights[43][24] = 16'sd-22;
        fc2_weights[43][25] = 16'sd1;
        fc2_weights[43][26] = 16'sd-17;
        fc2_weights[43][27] = 16'sd19;
        fc2_weights[43][28] = 16'sd-26;
        fc2_weights[43][29] = 16'sd-1;
        fc2_weights[43][30] = 16'sd5;
        fc2_weights[43][31] = 16'sd-21;
        fc2_weights[43][32] = 16'sd-10;
        fc2_weights[43][33] = 16'sd30;
        fc2_weights[43][34] = 16'sd-16;
        fc2_weights[43][35] = 16'sd4;
        fc2_weights[43][36] = 16'sd-24;
        fc2_weights[43][37] = 16'sd19;
        fc2_weights[43][38] = 16'sd-42;
        fc2_weights[43][39] = 16'sd-36;
        fc2_weights[43][40] = 16'sd56;
        fc2_weights[43][41] = 16'sd-41;
        fc2_weights[43][42] = 16'sd-27;
        fc2_weights[43][43] = 16'sd-32;
        fc2_weights[43][44] = 16'sd-23;
        fc2_weights[43][45] = 16'sd35;
        fc2_weights[43][46] = 16'sd-75;
        fc2_weights[43][47] = 16'sd-15;
        fc2_weights[43][48] = 16'sd-14;
        fc2_weights[43][49] = 16'sd-26;
        fc2_weights[43][50] = 16'sd-29;
        fc2_weights[43][51] = 16'sd30;
        fc2_weights[43][52] = 16'sd29;
        fc2_weights[43][53] = 16'sd-10;
        fc2_weights[43][54] = 16'sd-22;
        fc2_weights[43][55] = 16'sd18;
        fc2_weights[43][56] = 16'sd-13;
        fc2_weights[43][57] = 16'sd0;
        fc2_weights[43][58] = 16'sd19;
        fc2_weights[43][59] = 16'sd-48;
        fc2_weights[43][60] = 16'sd16;
        fc2_weights[43][61] = 16'sd93;
        fc2_weights[43][62] = 16'sd-21;
        fc2_weights[43][63] = 16'sd5;
        fc2_weights[43][64] = 16'sd-21;
        fc2_weights[43][65] = 16'sd2;
        fc2_weights[43][66] = 16'sd33;
        fc2_weights[43][67] = 16'sd14;
        fc2_weights[43][68] = 16'sd-4;
        fc2_weights[43][69] = 16'sd50;
        fc2_weights[43][70] = 16'sd-39;
        fc2_weights[43][71] = 16'sd5;
        fc2_weights[43][72] = 16'sd-29;
        fc2_weights[43][73] = 16'sd-53;
        fc2_weights[43][74] = 16'sd-13;
        fc2_weights[43][75] = 16'sd26;
        fc2_weights[43][76] = 16'sd29;
        fc2_weights[43][77] = 16'sd-36;
        fc2_weights[43][78] = 16'sd4;
        fc2_weights[43][79] = 16'sd-25;
        fc2_weights[43][80] = 16'sd-48;
        fc2_weights[43][81] = 16'sd12;
        fc2_weights[43][82] = 16'sd-15;
        fc2_weights[43][83] = 16'sd15;
        fc2_weights[43][84] = 16'sd-31;
        fc2_weights[43][85] = 16'sd35;
        fc2_weights[43][86] = 16'sd-46;
        fc2_weights[43][87] = 16'sd6;
        fc2_weights[43][88] = 16'sd-2;
        fc2_weights[43][89] = 16'sd38;
        fc2_weights[43][90] = 16'sd-33;
        fc2_weights[43][91] = 16'sd36;
        fc2_weights[43][92] = 16'sd-18;
        fc2_weights[43][93] = 16'sd-37;
        fc2_weights[43][94] = 16'sd-33;
        fc2_weights[43][95] = 16'sd21;
        fc2_weights[43][96] = 16'sd17;
        fc2_weights[43][97] = 16'sd-14;
        fc2_weights[43][98] = 16'sd7;
        fc2_weights[43][99] = 16'sd17;
        fc2_weights[43][100] = 16'sd9;
        fc2_weights[43][101] = 16'sd-31;
        fc2_weights[43][102] = 16'sd-21;
        fc2_weights[43][103] = 16'sd17;
        fc2_weights[43][104] = 16'sd-62;
        fc2_weights[43][105] = 16'sd34;
        fc2_weights[43][106] = 16'sd-17;
        fc2_weights[43][107] = 16'sd-24;
        fc2_weights[43][108] = 16'sd-30;
        fc2_weights[43][109] = 16'sd-49;
        fc2_weights[43][110] = 16'sd35;
        fc2_weights[43][111] = 16'sd-62;
        fc2_weights[43][112] = 16'sd5;
        fc2_weights[43][113] = 16'sd5;
        fc2_weights[43][114] = 16'sd1;
        fc2_weights[43][115] = 16'sd-2;
        fc2_weights[43][116] = 16'sd12;
        fc2_weights[43][117] = 16'sd22;
        fc2_weights[43][118] = 16'sd-41;
        fc2_weights[43][119] = 16'sd45;
        fc2_weights[43][120] = 16'sd-16;
        fc2_weights[43][121] = 16'sd-26;
        fc2_weights[43][122] = 16'sd26;
        fc2_weights[43][123] = 16'sd16;
        fc2_weights[43][124] = 16'sd-16;
        fc2_weights[43][125] = 16'sd15;
        fc2_weights[43][126] = 16'sd-18;
        fc2_weights[43][127] = 16'sd71;
        fc2_weights[44][0] = 16'sd-29;
        fc2_weights[44][1] = 16'sd-29;
        fc2_weights[44][2] = 16'sd21;
        fc2_weights[44][3] = 16'sd29;
        fc2_weights[44][4] = 16'sd-15;
        fc2_weights[44][5] = 16'sd-1;
        fc2_weights[44][6] = 16'sd-36;
        fc2_weights[44][7] = 16'sd-4;
        fc2_weights[44][8] = 16'sd-15;
        fc2_weights[44][9] = 16'sd7;
        fc2_weights[44][10] = 16'sd-28;
        fc2_weights[44][11] = 16'sd-23;
        fc2_weights[44][12] = 16'sd1;
        fc2_weights[44][13] = 16'sd48;
        fc2_weights[44][14] = 16'sd-2;
        fc2_weights[44][15] = 16'sd19;
        fc2_weights[44][16] = 16'sd-2;
        fc2_weights[44][17] = 16'sd15;
        fc2_weights[44][18] = 16'sd-28;
        fc2_weights[44][19] = 16'sd12;
        fc2_weights[44][20] = 16'sd4;
        fc2_weights[44][21] = 16'sd-11;
        fc2_weights[44][22] = 16'sd-10;
        fc2_weights[44][23] = 16'sd-31;
        fc2_weights[44][24] = 16'sd-36;
        fc2_weights[44][25] = 16'sd-1;
        fc2_weights[44][26] = 16'sd-10;
        fc2_weights[44][27] = 16'sd-1;
        fc2_weights[44][28] = 16'sd-11;
        fc2_weights[44][29] = 16'sd-37;
        fc2_weights[44][30] = 16'sd22;
        fc2_weights[44][31] = 16'sd-10;
        fc2_weights[44][32] = 16'sd15;
        fc2_weights[44][33] = 16'sd-7;
        fc2_weights[44][34] = 16'sd-6;
        fc2_weights[44][35] = 16'sd11;
        fc2_weights[44][36] = 16'sd-37;
        fc2_weights[44][37] = 16'sd-24;
        fc2_weights[44][38] = 16'sd-13;
        fc2_weights[44][39] = 16'sd-4;
        fc2_weights[44][40] = 16'sd33;
        fc2_weights[44][41] = 16'sd-31;
        fc2_weights[44][42] = 16'sd8;
        fc2_weights[44][43] = 16'sd-6;
        fc2_weights[44][44] = 16'sd32;
        fc2_weights[44][45] = 16'sd-4;
        fc2_weights[44][46] = 16'sd-27;
        fc2_weights[44][47] = 16'sd0;
        fc2_weights[44][48] = 16'sd8;
        fc2_weights[44][49] = 16'sd-1;
        fc2_weights[44][50] = 16'sd26;
        fc2_weights[44][51] = 16'sd-4;
        fc2_weights[44][52] = 16'sd1;
        fc2_weights[44][53] = 16'sd-11;
        fc2_weights[44][54] = 16'sd-46;
        fc2_weights[44][55] = 16'sd-8;
        fc2_weights[44][56] = 16'sd63;
        fc2_weights[44][57] = 16'sd34;
        fc2_weights[44][58] = 16'sd15;
        fc2_weights[44][59] = 16'sd-18;
        fc2_weights[44][60] = 16'sd-15;
        fc2_weights[44][61] = 16'sd-34;
        fc2_weights[44][62] = 16'sd-3;
        fc2_weights[44][63] = 16'sd-1;
        fc2_weights[44][64] = 16'sd-1;
        fc2_weights[44][65] = 16'sd14;
        fc2_weights[44][66] = 16'sd-22;
        fc2_weights[44][67] = 16'sd-15;
        fc2_weights[44][68] = 16'sd-17;
        fc2_weights[44][69] = 16'sd-11;
        fc2_weights[44][70] = 16'sd-28;
        fc2_weights[44][71] = 16'sd-5;
        fc2_weights[44][72] = 16'sd-21;
        fc2_weights[44][73] = 16'sd-26;
        fc2_weights[44][74] = 16'sd-6;
        fc2_weights[44][75] = 16'sd7;
        fc2_weights[44][76] = 16'sd-3;
        fc2_weights[44][77] = 16'sd-10;
        fc2_weights[44][78] = 16'sd17;
        fc2_weights[44][79] = 16'sd-1;
        fc2_weights[44][80] = 16'sd-22;
        fc2_weights[44][81] = 16'sd-19;
        fc2_weights[44][82] = 16'sd-35;
        fc2_weights[44][83] = 16'sd-25;
        fc2_weights[44][84] = 16'sd-21;
        fc2_weights[44][85] = 16'sd-4;
        fc2_weights[44][86] = 16'sd-16;
        fc2_weights[44][87] = 16'sd-7;
        fc2_weights[44][88] = 16'sd16;
        fc2_weights[44][89] = 16'sd-38;
        fc2_weights[44][90] = 16'sd-15;
        fc2_weights[44][91] = 16'sd8;
        fc2_weights[44][92] = 16'sd32;
        fc2_weights[44][93] = 16'sd-39;
        fc2_weights[44][94] = 16'sd7;
        fc2_weights[44][95] = 16'sd-35;
        fc2_weights[44][96] = 16'sd10;
        fc2_weights[44][97] = 16'sd-26;
        fc2_weights[44][98] = 16'sd-26;
        fc2_weights[44][99] = 16'sd-39;
        fc2_weights[44][100] = 16'sd27;
        fc2_weights[44][101] = 16'sd-26;
        fc2_weights[44][102] = 16'sd-2;
        fc2_weights[44][103] = 16'sd44;
        fc2_weights[44][104] = 16'sd43;
        fc2_weights[44][105] = 16'sd-26;
        fc2_weights[44][106] = 16'sd-8;
        fc2_weights[44][107] = 16'sd17;
        fc2_weights[44][108] = 16'sd-21;
        fc2_weights[44][109] = 16'sd11;
        fc2_weights[44][110] = 16'sd62;
        fc2_weights[44][111] = 16'sd-20;
        fc2_weights[44][112] = 16'sd-12;
        fc2_weights[44][113] = 16'sd-40;
        fc2_weights[44][114] = 16'sd-1;
        fc2_weights[44][115] = 16'sd-20;
        fc2_weights[44][116] = 16'sd-15;
        fc2_weights[44][117] = 16'sd-21;
        fc2_weights[44][118] = 16'sd-43;
        fc2_weights[44][119] = 16'sd-37;
        fc2_weights[44][120] = 16'sd-21;
        fc2_weights[44][121] = 16'sd-23;
        fc2_weights[44][122] = 16'sd-32;
        fc2_weights[44][123] = 16'sd37;
        fc2_weights[44][124] = 16'sd-24;
        fc2_weights[44][125] = 16'sd-7;
        fc2_weights[44][126] = 16'sd21;
        fc2_weights[44][127] = 16'sd-53;
        fc2_weights[45][0] = 16'sd18;
        fc2_weights[45][1] = 16'sd-3;
        fc2_weights[45][2] = 16'sd16;
        fc2_weights[45][3] = 16'sd39;
        fc2_weights[45][4] = 16'sd37;
        fc2_weights[45][5] = 16'sd10;
        fc2_weights[45][6] = 16'sd-43;
        fc2_weights[45][7] = 16'sd-8;
        fc2_weights[45][8] = 16'sd-70;
        fc2_weights[45][9] = 16'sd-5;
        fc2_weights[45][10] = 16'sd7;
        fc2_weights[45][11] = 16'sd-32;
        fc2_weights[45][12] = 16'sd-16;
        fc2_weights[45][13] = 16'sd3;
        fc2_weights[45][14] = 16'sd0;
        fc2_weights[45][15] = 16'sd44;
        fc2_weights[45][16] = 16'sd22;
        fc2_weights[45][17] = 16'sd24;
        fc2_weights[45][18] = 16'sd1;
        fc2_weights[45][19] = 16'sd25;
        fc2_weights[45][20] = 16'sd-14;
        fc2_weights[45][21] = 16'sd-44;
        fc2_weights[45][22] = 16'sd-40;
        fc2_weights[45][23] = 16'sd-13;
        fc2_weights[45][24] = 16'sd-4;
        fc2_weights[45][25] = 16'sd-5;
        fc2_weights[45][26] = 16'sd-14;
        fc2_weights[45][27] = 16'sd20;
        fc2_weights[45][28] = 16'sd-4;
        fc2_weights[45][29] = 16'sd-36;
        fc2_weights[45][30] = 16'sd-17;
        fc2_weights[45][31] = 16'sd-19;
        fc2_weights[45][32] = 16'sd-45;
        fc2_weights[45][33] = 16'sd-40;
        fc2_weights[45][34] = 16'sd43;
        fc2_weights[45][35] = 16'sd31;
        fc2_weights[45][36] = 16'sd-37;
        fc2_weights[45][37] = 16'sd-19;
        fc2_weights[45][38] = 16'sd17;
        fc2_weights[45][39] = 16'sd-19;
        fc2_weights[45][40] = 16'sd22;
        fc2_weights[45][41] = 16'sd-4;
        fc2_weights[45][42] = 16'sd-3;
        fc2_weights[45][43] = 16'sd-25;
        fc2_weights[45][44] = 16'sd47;
        fc2_weights[45][45] = 16'sd22;
        fc2_weights[45][46] = 16'sd53;
        fc2_weights[45][47] = 16'sd-14;
        fc2_weights[45][48] = 16'sd22;
        fc2_weights[45][49] = 16'sd-2;
        fc2_weights[45][50] = 16'sd-14;
        fc2_weights[45][51] = 16'sd-15;
        fc2_weights[45][52] = 16'sd-16;
        fc2_weights[45][53] = 16'sd-98;
        fc2_weights[45][54] = 16'sd-30;
        fc2_weights[45][55] = 16'sd-40;
        fc2_weights[45][56] = 16'sd26;
        fc2_weights[45][57] = 16'sd20;
        fc2_weights[45][58] = 16'sd0;
        fc2_weights[45][59] = 16'sd27;
        fc2_weights[45][60] = 16'sd-8;
        fc2_weights[45][61] = 16'sd-48;
        fc2_weights[45][62] = 16'sd16;
        fc2_weights[45][63] = 16'sd7;
        fc2_weights[45][64] = 16'sd-16;
        fc2_weights[45][65] = 16'sd44;
        fc2_weights[45][66] = 16'sd20;
        fc2_weights[45][67] = 16'sd-18;
        fc2_weights[45][68] = 16'sd8;
        fc2_weights[45][69] = 16'sd26;
        fc2_weights[45][70] = 16'sd-38;
        fc2_weights[45][71] = 16'sd33;
        fc2_weights[45][72] = 16'sd-20;
        fc2_weights[45][73] = 16'sd-12;
        fc2_weights[45][74] = 16'sd14;
        fc2_weights[45][75] = 16'sd-31;
        fc2_weights[45][76] = 16'sd-34;
        fc2_weights[45][77] = 16'sd9;
        fc2_weights[45][78] = 16'sd-14;
        fc2_weights[45][79] = 16'sd-40;
        fc2_weights[45][80] = 16'sd-13;
        fc2_weights[45][81] = 16'sd8;
        fc2_weights[45][82] = 16'sd-45;
        fc2_weights[45][83] = 16'sd-13;
        fc2_weights[45][84] = 16'sd0;
        fc2_weights[45][85] = 16'sd-20;
        fc2_weights[45][86] = 16'sd-30;
        fc2_weights[45][87] = 16'sd1;
        fc2_weights[45][88] = 16'sd-6;
        fc2_weights[45][89] = 16'sd18;
        fc2_weights[45][90] = 16'sd-3;
        fc2_weights[45][91] = 16'sd-19;
        fc2_weights[45][92] = 16'sd-17;
        fc2_weights[45][93] = 16'sd-37;
        fc2_weights[45][94] = 16'sd28;
        fc2_weights[45][95] = 16'sd-27;
        fc2_weights[45][96] = 16'sd48;
        fc2_weights[45][97] = 16'sd-10;
        fc2_weights[45][98] = 16'sd-2;
        fc2_weights[45][99] = 16'sd-24;
        fc2_weights[45][100] = 16'sd21;
        fc2_weights[45][101] = 16'sd19;
        fc2_weights[45][102] = 16'sd54;
        fc2_weights[45][103] = 16'sd-61;
        fc2_weights[45][104] = 16'sd126;
        fc2_weights[45][105] = 16'sd-7;
        fc2_weights[45][106] = 16'sd-10;
        fc2_weights[45][107] = 16'sd12;
        fc2_weights[45][108] = 16'sd-32;
        fc2_weights[45][109] = 16'sd-79;
        fc2_weights[45][110] = 16'sd46;
        fc2_weights[45][111] = 16'sd28;
        fc2_weights[45][112] = 16'sd-57;
        fc2_weights[45][113] = 16'sd-56;
        fc2_weights[45][114] = 16'sd49;
        fc2_weights[45][115] = 16'sd6;
        fc2_weights[45][116] = 16'sd-11;
        fc2_weights[45][117] = 16'sd-21;
        fc2_weights[45][118] = 16'sd-20;
        fc2_weights[45][119] = 16'sd-13;
        fc2_weights[45][120] = 16'sd-35;
        fc2_weights[45][121] = 16'sd-35;
        fc2_weights[45][122] = 16'sd-1;
        fc2_weights[45][123] = 16'sd88;
        fc2_weights[45][124] = 16'sd-25;
        fc2_weights[45][125] = 16'sd58;
        fc2_weights[45][126] = 16'sd-7;
        fc2_weights[45][127] = 16'sd-34;
        fc2_weights[46][0] = 16'sd76;
        fc2_weights[46][1] = 16'sd-20;
        fc2_weights[46][2] = 16'sd5;
        fc2_weights[46][3] = 16'sd-51;
        fc2_weights[46][4] = 16'sd15;
        fc2_weights[46][5] = 16'sd9;
        fc2_weights[46][6] = 16'sd45;
        fc2_weights[46][7] = 16'sd-59;
        fc2_weights[46][8] = 16'sd59;
        fc2_weights[46][9] = 16'sd33;
        fc2_weights[46][10] = 16'sd1;
        fc2_weights[46][11] = 16'sd-18;
        fc2_weights[46][12] = 16'sd42;
        fc2_weights[46][13] = 16'sd-37;
        fc2_weights[46][14] = 16'sd-19;
        fc2_weights[46][15] = 16'sd-13;
        fc2_weights[46][16] = 16'sd-22;
        fc2_weights[46][17] = 16'sd9;
        fc2_weights[46][18] = 16'sd51;
        fc2_weights[46][19] = 16'sd-58;
        fc2_weights[46][20] = 16'sd34;
        fc2_weights[46][21] = 16'sd7;
        fc2_weights[46][22] = 16'sd27;
        fc2_weights[46][23] = 16'sd27;
        fc2_weights[46][24] = 16'sd-56;
        fc2_weights[46][25] = 16'sd-33;
        fc2_weights[46][26] = 16'sd8;
        fc2_weights[46][27] = 16'sd1;
        fc2_weights[46][28] = 16'sd17;
        fc2_weights[46][29] = 16'sd-45;
        fc2_weights[46][30] = 16'sd23;
        fc2_weights[46][31] = 16'sd17;
        fc2_weights[46][32] = 16'sd-4;
        fc2_weights[46][33] = 16'sd38;
        fc2_weights[46][34] = 16'sd-42;
        fc2_weights[46][35] = 16'sd-25;
        fc2_weights[46][36] = 16'sd13;
        fc2_weights[46][37] = 16'sd15;
        fc2_weights[46][38] = 16'sd8;
        fc2_weights[46][39] = 16'sd30;
        fc2_weights[46][40] = 16'sd-43;
        fc2_weights[46][41] = 16'sd-51;
        fc2_weights[46][42] = 16'sd0;
        fc2_weights[46][43] = 16'sd44;
        fc2_weights[46][44] = 16'sd-83;
        fc2_weights[46][45] = 16'sd-76;
        fc2_weights[46][46] = 16'sd-56;
        fc2_weights[46][47] = 16'sd-9;
        fc2_weights[46][48] = 16'sd-1;
        fc2_weights[46][49] = 16'sd-42;
        fc2_weights[46][50] = 16'sd46;
        fc2_weights[46][51] = 16'sd-38;
        fc2_weights[46][52] = 16'sd-56;
        fc2_weights[46][53] = 16'sd46;
        fc2_weights[46][54] = 16'sd48;
        fc2_weights[46][55] = 16'sd-4;
        fc2_weights[46][56] = 16'sd-3;
        fc2_weights[46][57] = 16'sd-88;
        fc2_weights[46][58] = 16'sd9;
        fc2_weights[46][59] = 16'sd7;
        fc2_weights[46][60] = 16'sd-37;
        fc2_weights[46][61] = 16'sd-7;
        fc2_weights[46][62] = 16'sd-59;
        fc2_weights[46][63] = 16'sd-50;
        fc2_weights[46][64] = 16'sd-5;
        fc2_weights[46][65] = 16'sd-42;
        fc2_weights[46][66] = 16'sd-57;
        fc2_weights[46][67] = 16'sd-9;
        fc2_weights[46][68] = 16'sd20;
        fc2_weights[46][69] = 16'sd-37;
        fc2_weights[46][70] = 16'sd32;
        fc2_weights[46][71] = 16'sd10;
        fc2_weights[46][72] = 16'sd105;
        fc2_weights[46][73] = 16'sd12;
        fc2_weights[46][74] = 16'sd-73;
        fc2_weights[46][75] = 16'sd-8;
        fc2_weights[46][76] = 16'sd-47;
        fc2_weights[46][77] = 16'sd-18;
        fc2_weights[46][78] = 16'sd2;
        fc2_weights[46][79] = 16'sd-30;
        fc2_weights[46][80] = 16'sd17;
        fc2_weights[46][81] = 16'sd-36;
        fc2_weights[46][82] = 16'sd-2;
        fc2_weights[46][83] = 16'sd8;
        fc2_weights[46][84] = 16'sd-52;
        fc2_weights[46][85] = 16'sd-22;
        fc2_weights[46][86] = 16'sd-37;
        fc2_weights[46][87] = 16'sd-23;
        fc2_weights[46][88] = 16'sd16;
        fc2_weights[46][89] = 16'sd1;
        fc2_weights[46][90] = 16'sd-97;
        fc2_weights[46][91] = 16'sd-67;
        fc2_weights[46][92] = 16'sd-49;
        fc2_weights[46][93] = 16'sd20;
        fc2_weights[46][94] = 16'sd4;
        fc2_weights[46][95] = 16'sd-16;
        fc2_weights[46][96] = 16'sd-36;
        fc2_weights[46][97] = 16'sd81;
        fc2_weights[46][98] = 16'sd-34;
        fc2_weights[46][99] = 16'sd13;
        fc2_weights[46][100] = 16'sd-62;
        fc2_weights[46][101] = 16'sd-4;
        fc2_weights[46][102] = 16'sd16;
        fc2_weights[46][103] = 16'sd-70;
        fc2_weights[46][104] = 16'sd-78;
        fc2_weights[46][105] = 16'sd41;
        fc2_weights[46][106] = 16'sd16;
        fc2_weights[46][107] = 16'sd-26;
        fc2_weights[46][108] = 16'sd46;
        fc2_weights[46][109] = 16'sd31;
        fc2_weights[46][110] = 16'sd-36;
        fc2_weights[46][111] = 16'sd-75;
        fc2_weights[46][112] = 16'sd50;
        fc2_weights[46][113] = 16'sd26;
        fc2_weights[46][114] = 16'sd30;
        fc2_weights[46][115] = 16'sd24;
        fc2_weights[46][116] = 16'sd-17;
        fc2_weights[46][117] = 16'sd14;
        fc2_weights[46][118] = 16'sd100;
        fc2_weights[46][119] = 16'sd-35;
        fc2_weights[46][120] = 16'sd23;
        fc2_weights[46][121] = 16'sd20;
        fc2_weights[46][122] = 16'sd-13;
        fc2_weights[46][123] = 16'sd-79;
        fc2_weights[46][124] = 16'sd67;
        fc2_weights[46][125] = 16'sd-76;
        fc2_weights[46][126] = 16'sd-89;
        fc2_weights[46][127] = 16'sd-6;
        fc2_weights[47][0] = 16'sd-70;
        fc2_weights[47][1] = 16'sd16;
        fc2_weights[47][2] = 16'sd-43;
        fc2_weights[47][3] = 16'sd-40;
        fc2_weights[47][4] = 16'sd31;
        fc2_weights[47][5] = 16'sd0;
        fc2_weights[47][6] = 16'sd-17;
        fc2_weights[47][7] = 16'sd13;
        fc2_weights[47][8] = 16'sd50;
        fc2_weights[47][9] = 16'sd-32;
        fc2_weights[47][10] = 16'sd-21;
        fc2_weights[47][11] = 16'sd50;
        fc2_weights[47][12] = 16'sd21;
        fc2_weights[47][13] = 16'sd9;
        fc2_weights[47][14] = 16'sd-43;
        fc2_weights[47][15] = 16'sd-23;
        fc2_weights[47][16] = 16'sd-47;
        fc2_weights[47][17] = 16'sd9;
        fc2_weights[47][18] = 16'sd-7;
        fc2_weights[47][19] = 16'sd-45;
        fc2_weights[47][20] = 16'sd19;
        fc2_weights[47][21] = 16'sd20;
        fc2_weights[47][22] = 16'sd61;
        fc2_weights[47][23] = 16'sd-2;
        fc2_weights[47][24] = 16'sd-30;
        fc2_weights[47][25] = 16'sd37;
        fc2_weights[47][26] = 16'sd19;
        fc2_weights[47][27] = 16'sd-27;
        fc2_weights[47][28] = 16'sd-26;
        fc2_weights[47][29] = 16'sd13;
        fc2_weights[47][30] = 16'sd-10;
        fc2_weights[47][31] = 16'sd-10;
        fc2_weights[47][32] = 16'sd-57;
        fc2_weights[47][33] = 16'sd2;
        fc2_weights[47][34] = 16'sd-13;
        fc2_weights[47][35] = 16'sd-80;
        fc2_weights[47][36] = 16'sd2;
        fc2_weights[47][37] = 16'sd-10;
        fc2_weights[47][38] = 16'sd27;
        fc2_weights[47][39] = 16'sd36;
        fc2_weights[47][40] = 16'sd-4;
        fc2_weights[47][41] = 16'sd-16;
        fc2_weights[47][42] = 16'sd58;
        fc2_weights[47][43] = 16'sd-8;
        fc2_weights[47][44] = 16'sd-15;
        fc2_weights[47][45] = 16'sd-30;
        fc2_weights[47][46] = 16'sd-49;
        fc2_weights[47][47] = 16'sd-19;
        fc2_weights[47][48] = 16'sd-36;
        fc2_weights[47][49] = 16'sd7;
        fc2_weights[47][50] = 16'sd-30;
        fc2_weights[47][51] = 16'sd-66;
        fc2_weights[47][52] = 16'sd-51;
        fc2_weights[47][53] = 16'sd-20;
        fc2_weights[47][54] = 16'sd-5;
        fc2_weights[47][55] = 16'sd-57;
        fc2_weights[47][56] = 16'sd0;
        fc2_weights[47][57] = 16'sd-52;
        fc2_weights[47][58] = 16'sd-26;
        fc2_weights[47][59] = 16'sd-21;
        fc2_weights[47][60] = 16'sd2;
        fc2_weights[47][61] = 16'sd28;
        fc2_weights[47][62] = 16'sd-54;
        fc2_weights[47][63] = 16'sd-31;
        fc2_weights[47][64] = 16'sd-56;
        fc2_weights[47][65] = 16'sd-67;
        fc2_weights[47][66] = 16'sd-27;
        fc2_weights[47][67] = 16'sd-28;
        fc2_weights[47][68] = 16'sd26;
        fc2_weights[47][69] = 16'sd-56;
        fc2_weights[47][70] = 16'sd8;
        fc2_weights[47][71] = 16'sd-65;
        fc2_weights[47][72] = 16'sd-31;
        fc2_weights[47][73] = 16'sd31;
        fc2_weights[47][74] = 16'sd-10;
        fc2_weights[47][75] = 16'sd-23;
        fc2_weights[47][76] = 16'sd35;
        fc2_weights[47][77] = 16'sd-38;
        fc2_weights[47][78] = 16'sd31;
        fc2_weights[47][79] = 16'sd23;
        fc2_weights[47][80] = 16'sd-43;
        fc2_weights[47][81] = 16'sd-55;
        fc2_weights[47][82] = 16'sd13;
        fc2_weights[47][83] = 16'sd-21;
        fc2_weights[47][84] = 16'sd-41;
        fc2_weights[47][85] = 16'sd-22;
        fc2_weights[47][86] = 16'sd-45;
        fc2_weights[47][87] = 16'sd22;
        fc2_weights[47][88] = 16'sd19;
        fc2_weights[47][89] = 16'sd32;
        fc2_weights[47][90] = 16'sd-28;
        fc2_weights[47][91] = 16'sd-38;
        fc2_weights[47][92] = 16'sd-1;
        fc2_weights[47][93] = 16'sd-51;
        fc2_weights[47][94] = 16'sd-56;
        fc2_weights[47][95] = 16'sd32;
        fc2_weights[47][96] = 16'sd-44;
        fc2_weights[47][97] = 16'sd11;
        fc2_weights[47][98] = 16'sd-51;
        fc2_weights[47][99] = 16'sd-5;
        fc2_weights[47][100] = 16'sd-23;
        fc2_weights[47][101] = 16'sd-15;
        fc2_weights[47][102] = 16'sd-36;
        fc2_weights[47][103] = 16'sd-78;
        fc2_weights[47][104] = 16'sd-33;
        fc2_weights[47][105] = 16'sd-36;
        fc2_weights[47][106] = 16'sd-1;
        fc2_weights[47][107] = 16'sd7;
        fc2_weights[47][108] = 16'sd7;
        fc2_weights[47][109] = 16'sd-43;
        fc2_weights[47][110] = 16'sd-16;
        fc2_weights[47][111] = 16'sd8;
        fc2_weights[47][112] = 16'sd7;
        fc2_weights[47][113] = 16'sd88;
        fc2_weights[47][114] = 16'sd3;
        fc2_weights[47][115] = 16'sd-3;
        fc2_weights[47][116] = 16'sd6;
        fc2_weights[47][117] = 16'sd-34;
        fc2_weights[47][118] = 16'sd54;
        fc2_weights[47][119] = 16'sd1;
        fc2_weights[47][120] = 16'sd41;
        fc2_weights[47][121] = 16'sd13;
        fc2_weights[47][122] = 16'sd-33;
        fc2_weights[47][123] = 16'sd-88;
        fc2_weights[47][124] = 16'sd42;
        fc2_weights[47][125] = 16'sd-41;
        fc2_weights[47][126] = 16'sd-74;
        fc2_weights[47][127] = 16'sd-3;
        fc2_weights[48][0] = 16'sd-1;
        fc2_weights[48][1] = 16'sd-48;
        fc2_weights[48][2] = 16'sd1;
        fc2_weights[48][3] = 16'sd-9;
        fc2_weights[48][4] = 16'sd-13;
        fc2_weights[48][5] = 16'sd-56;
        fc2_weights[48][6] = 16'sd-71;
        fc2_weights[48][7] = 16'sd-70;
        fc2_weights[48][8] = 16'sd-44;
        fc2_weights[48][9] = 16'sd-32;
        fc2_weights[48][10] = 16'sd-38;
        fc2_weights[48][11] = 16'sd-32;
        fc2_weights[48][12] = 16'sd-45;
        fc2_weights[48][13] = 16'sd7;
        fc2_weights[48][14] = 16'sd76;
        fc2_weights[48][15] = 16'sd3;
        fc2_weights[48][16] = 16'sd34;
        fc2_weights[48][17] = 16'sd-23;
        fc2_weights[48][18] = 16'sd8;
        fc2_weights[48][19] = 16'sd4;
        fc2_weights[48][20] = 16'sd11;
        fc2_weights[48][21] = 16'sd-57;
        fc2_weights[48][22] = 16'sd-70;
        fc2_weights[48][23] = 16'sd-40;
        fc2_weights[48][24] = 16'sd31;
        fc2_weights[48][25] = 16'sd69;
        fc2_weights[48][26] = 16'sd-65;
        fc2_weights[48][27] = 16'sd12;
        fc2_weights[48][28] = 16'sd-16;
        fc2_weights[48][29] = 16'sd-51;
        fc2_weights[48][30] = 16'sd15;
        fc2_weights[48][31] = 16'sd-70;
        fc2_weights[48][32] = 16'sd-75;
        fc2_weights[48][33] = 16'sd-37;
        fc2_weights[48][34] = 16'sd11;
        fc2_weights[48][35] = 16'sd30;
        fc2_weights[48][36] = 16'sd-81;
        fc2_weights[48][37] = 16'sd-74;
        fc2_weights[48][38] = 16'sd10;
        fc2_weights[48][39] = 16'sd16;
        fc2_weights[48][40] = 16'sd-26;
        fc2_weights[48][41] = 16'sd-16;
        fc2_weights[48][42] = 16'sd-7;
        fc2_weights[48][43] = 16'sd-9;
        fc2_weights[48][44] = 16'sd81;
        fc2_weights[48][45] = 16'sd42;
        fc2_weights[48][46] = 16'sd38;
        fc2_weights[48][47] = 16'sd-24;
        fc2_weights[48][48] = 16'sd15;
        fc2_weights[48][49] = 16'sd16;
        fc2_weights[48][50] = 16'sd30;
        fc2_weights[48][51] = 16'sd-5;
        fc2_weights[48][52] = 16'sd8;
        fc2_weights[48][53] = 16'sd14;
        fc2_weights[48][54] = 16'sd-91;
        fc2_weights[48][55] = 16'sd-52;
        fc2_weights[48][56] = 16'sd48;
        fc2_weights[48][57] = 16'sd38;
        fc2_weights[48][58] = 16'sd34;
        fc2_weights[48][59] = 16'sd29;
        fc2_weights[48][60] = 16'sd-26;
        fc2_weights[48][61] = 16'sd-90;
        fc2_weights[48][62] = 16'sd37;
        fc2_weights[48][63] = 16'sd25;
        fc2_weights[48][64] = 16'sd-53;
        fc2_weights[48][65] = 16'sd76;
        fc2_weights[48][66] = 16'sd44;
        fc2_weights[48][67] = 16'sd-24;
        fc2_weights[48][68] = 16'sd0;
        fc2_weights[48][69] = 16'sd52;
        fc2_weights[48][70] = 16'sd-10;
        fc2_weights[48][71] = 16'sd13;
        fc2_weights[48][72] = 16'sd-6;
        fc2_weights[48][73] = 16'sd-31;
        fc2_weights[48][74] = 16'sd41;
        fc2_weights[48][75] = 16'sd-8;
        fc2_weights[48][76] = 16'sd-18;
        fc2_weights[48][77] = 16'sd26;
        fc2_weights[48][78] = 16'sd-1;
        fc2_weights[48][79] = 16'sd-27;
        fc2_weights[48][80] = 16'sd-47;
        fc2_weights[48][81] = 16'sd33;
        fc2_weights[48][82] = 16'sd-44;
        fc2_weights[48][83] = 16'sd4;
        fc2_weights[48][84] = 16'sd-26;
        fc2_weights[48][85] = 16'sd-36;
        fc2_weights[48][86] = 16'sd-26;
        fc2_weights[48][87] = 16'sd-6;
        fc2_weights[48][88] = 16'sd67;
        fc2_weights[48][89] = 16'sd13;
        fc2_weights[48][90] = 16'sd53;
        fc2_weights[48][91] = 16'sd-41;
        fc2_weights[48][92] = 16'sd0;
        fc2_weights[48][93] = 16'sd-61;
        fc2_weights[48][94] = 16'sd-10;
        fc2_weights[48][95] = 16'sd-66;
        fc2_weights[48][96] = 16'sd113;
        fc2_weights[48][97] = 16'sd5;
        fc2_weights[48][98] = 16'sd75;
        fc2_weights[48][99] = 16'sd-25;
        fc2_weights[48][100] = 16'sd24;
        fc2_weights[48][101] = 16'sd-6;
        fc2_weights[48][102] = 16'sd53;
        fc2_weights[48][103] = 16'sd-59;
        fc2_weights[48][104] = 16'sd39;
        fc2_weights[48][105] = 16'sd-21;
        fc2_weights[48][106] = 16'sd10;
        fc2_weights[48][107] = 16'sd59;
        fc2_weights[48][108] = 16'sd-31;
        fc2_weights[48][109] = 16'sd-12;
        fc2_weights[48][110] = 16'sd82;
        fc2_weights[48][111] = 16'sd8;
        fc2_weights[48][112] = 16'sd-41;
        fc2_weights[48][113] = 16'sd-81;
        fc2_weights[48][114] = 16'sd-1;
        fc2_weights[48][115] = 16'sd-64;
        fc2_weights[48][116] = 16'sd2;
        fc2_weights[48][117] = 16'sd-14;
        fc2_weights[48][118] = 16'sd24;
        fc2_weights[48][119] = 16'sd-48;
        fc2_weights[48][120] = 16'sd-29;
        fc2_weights[48][121] = 16'sd53;
        fc2_weights[48][122] = 16'sd9;
        fc2_weights[48][123] = 16'sd105;
        fc2_weights[48][124] = 16'sd-5;
        fc2_weights[48][125] = 16'sd-12;
        fc2_weights[48][126] = 16'sd12;
        fc2_weights[48][127] = 16'sd-67;
        fc2_weights[49][0] = 16'sd-3;
        fc2_weights[49][1] = 16'sd-73;
        fc2_weights[49][2] = 16'sd-44;
        fc2_weights[49][3] = 16'sd-52;
        fc2_weights[49][4] = 16'sd28;
        fc2_weights[49][5] = 16'sd18;
        fc2_weights[49][6] = 16'sd-22;
        fc2_weights[49][7] = 16'sd25;
        fc2_weights[49][8] = 16'sd4;
        fc2_weights[49][9] = 16'sd-56;
        fc2_weights[49][10] = 16'sd36;
        fc2_weights[49][11] = 16'sd39;
        fc2_weights[49][12] = 16'sd-31;
        fc2_weights[49][13] = 16'sd-74;
        fc2_weights[49][14] = 16'sd14;
        fc2_weights[49][15] = 16'sd-38;
        fc2_weights[49][16] = 16'sd47;
        fc2_weights[49][17] = 16'sd-29;
        fc2_weights[49][18] = 16'sd-24;
        fc2_weights[49][19] = 16'sd-3;
        fc2_weights[49][20] = 16'sd-51;
        fc2_weights[49][21] = 16'sd-17;
        fc2_weights[49][22] = 16'sd39;
        fc2_weights[49][23] = 16'sd32;
        fc2_weights[49][24] = 16'sd-5;
        fc2_weights[49][25] = 16'sd45;
        fc2_weights[49][26] = 16'sd38;
        fc2_weights[49][27] = 16'sd-31;
        fc2_weights[49][28] = 16'sd14;
        fc2_weights[49][29] = 16'sd78;
        fc2_weights[49][30] = 16'sd-15;
        fc2_weights[49][31] = 16'sd8;
        fc2_weights[49][32] = 16'sd-41;
        fc2_weights[49][33] = 16'sd5;
        fc2_weights[49][34] = 16'sd-56;
        fc2_weights[49][35] = 16'sd30;
        fc2_weights[49][36] = 16'sd13;
        fc2_weights[49][37] = 16'sd-95;
        fc2_weights[49][38] = 16'sd33;
        fc2_weights[49][39] = 16'sd54;
        fc2_weights[49][40] = 16'sd-71;
        fc2_weights[49][41] = 16'sd92;
        fc2_weights[49][42] = 16'sd11;
        fc2_weights[49][43] = 16'sd-43;
        fc2_weights[49][44] = 16'sd4;
        fc2_weights[49][45] = 16'sd26;
        fc2_weights[49][46] = 16'sd52;
        fc2_weights[49][47] = 16'sd12;
        fc2_weights[49][48] = 16'sd-38;
        fc2_weights[49][49] = 16'sd66;
        fc2_weights[49][50] = 16'sd-7;
        fc2_weights[49][51] = 16'sd63;
        fc2_weights[49][52] = 16'sd-47;
        fc2_weights[49][53] = 16'sd-18;
        fc2_weights[49][54] = 16'sd51;
        fc2_weights[49][55] = 16'sd49;
        fc2_weights[49][56] = 16'sd19;
        fc2_weights[49][57] = 16'sd6;
        fc2_weights[49][58] = 16'sd-49;
        fc2_weights[49][59] = 16'sd-21;
        fc2_weights[49][60] = 16'sd46;
        fc2_weights[49][61] = 16'sd-12;
        fc2_weights[49][62] = 16'sd41;
        fc2_weights[49][63] = 16'sd-44;
        fc2_weights[49][64] = 16'sd41;
        fc2_weights[49][65] = 16'sd27;
        fc2_weights[49][66] = 16'sd12;
        fc2_weights[49][67] = 16'sd19;
        fc2_weights[49][68] = 16'sd-57;
        fc2_weights[49][69] = 16'sd-42;
        fc2_weights[49][70] = 16'sd-11;
        fc2_weights[49][71] = 16'sd51;
        fc2_weights[49][72] = 16'sd-47;
        fc2_weights[49][73] = 16'sd-24;
        fc2_weights[49][74] = 16'sd-31;
        fc2_weights[49][75] = 16'sd-7;
        fc2_weights[49][76] = 16'sd19;
        fc2_weights[49][77] = 16'sd118;
        fc2_weights[49][78] = 16'sd-19;
        fc2_weights[49][79] = 16'sd11;
        fc2_weights[49][80] = 16'sd-10;
        fc2_weights[49][81] = 16'sd1;
        fc2_weights[49][82] = 16'sd42;
        fc2_weights[49][83] = 16'sd31;
        fc2_weights[49][84] = 16'sd-26;
        fc2_weights[49][85] = 16'sd-8;
        fc2_weights[49][86] = 16'sd7;
        fc2_weights[49][87] = 16'sd-93;
        fc2_weights[49][88] = 16'sd26;
        fc2_weights[49][89] = 16'sd28;
        fc2_weights[49][90] = 16'sd-12;
        fc2_weights[49][91] = 16'sd12;
        fc2_weights[49][92] = 16'sd11;
        fc2_weights[49][93] = 16'sd7;
        fc2_weights[49][94] = 16'sd-71;
        fc2_weights[49][95] = 16'sd41;
        fc2_weights[49][96] = 16'sd-2;
        fc2_weights[49][97] = 16'sd73;
        fc2_weights[49][98] = 16'sd86;
        fc2_weights[49][99] = 16'sd46;
        fc2_weights[49][100] = 16'sd43;
        fc2_weights[49][101] = 16'sd-10;
        fc2_weights[49][102] = 16'sd-39;
        fc2_weights[49][103] = 16'sd-18;
        fc2_weights[49][104] = 16'sd49;
        fc2_weights[49][105] = 16'sd-26;
        fc2_weights[49][106] = 16'sd-8;
        fc2_weights[49][107] = 16'sd60;
        fc2_weights[49][108] = 16'sd-54;
        fc2_weights[49][109] = 16'sd19;
        fc2_weights[49][110] = 16'sd-3;
        fc2_weights[49][111] = 16'sd39;
        fc2_weights[49][112] = 16'sd-32;
        fc2_weights[49][113] = 16'sd7;
        fc2_weights[49][114] = 16'sd28;
        fc2_weights[49][115] = 16'sd28;
        fc2_weights[49][116] = 16'sd-24;
        fc2_weights[49][117] = 16'sd-6;
        fc2_weights[49][118] = 16'sd32;
        fc2_weights[49][119] = 16'sd-17;
        fc2_weights[49][120] = 16'sd-55;
        fc2_weights[49][121] = 16'sd58;
        fc2_weights[49][122] = 16'sd57;
        fc2_weights[49][123] = 16'sd21;
        fc2_weights[49][124] = 16'sd0;
        fc2_weights[49][125] = 16'sd-15;
        fc2_weights[49][126] = 16'sd25;
        fc2_weights[49][127] = 16'sd-17;
        fc2_weights[50][0] = 16'sd-14;
        fc2_weights[50][1] = 16'sd8;
        fc2_weights[50][2] = 16'sd-2;
        fc2_weights[50][3] = 16'sd84;
        fc2_weights[50][4] = 16'sd-50;
        fc2_weights[50][5] = 16'sd-23;
        fc2_weights[50][6] = 16'sd-14;
        fc2_weights[50][7] = 16'sd52;
        fc2_weights[50][8] = 16'sd109;
        fc2_weights[50][9] = 16'sd-18;
        fc2_weights[50][10] = 16'sd-46;
        fc2_weights[50][11] = 16'sd-51;
        fc2_weights[50][12] = 16'sd66;
        fc2_weights[50][13] = 16'sd4;
        fc2_weights[50][14] = 16'sd-34;
        fc2_weights[50][15] = 16'sd-24;
        fc2_weights[50][16] = 16'sd-31;
        fc2_weights[50][17] = 16'sd52;
        fc2_weights[50][18] = 16'sd2;
        fc2_weights[50][19] = 16'sd34;
        fc2_weights[50][20] = 16'sd-1;
        fc2_weights[50][21] = 16'sd15;
        fc2_weights[50][22] = 16'sd4;
        fc2_weights[50][23] = 16'sd-29;
        fc2_weights[50][24] = 16'sd-21;
        fc2_weights[50][25] = 16'sd-43;
        fc2_weights[50][26] = 16'sd16;
        fc2_weights[50][27] = 16'sd-45;
        fc2_weights[50][28] = 16'sd48;
        fc2_weights[50][29] = 16'sd11;
        fc2_weights[50][30] = 16'sd24;
        fc2_weights[50][31] = 16'sd48;
        fc2_weights[50][32] = 16'sd33;
        fc2_weights[50][33] = 16'sd30;
        fc2_weights[50][34] = 16'sd-7;
        fc2_weights[50][35] = 16'sd-26;
        fc2_weights[50][36] = 16'sd-32;
        fc2_weights[50][37] = 16'sd-15;
        fc2_weights[50][38] = 16'sd7;
        fc2_weights[50][39] = 16'sd-4;
        fc2_weights[50][40] = 16'sd47;
        fc2_weights[50][41] = 16'sd-51;
        fc2_weights[50][42] = 16'sd9;
        fc2_weights[50][43] = 16'sd62;
        fc2_weights[50][44] = 16'sd-16;
        fc2_weights[50][45] = 16'sd-48;
        fc2_weights[50][46] = 16'sd-66;
        fc2_weights[50][47] = 16'sd2;
        fc2_weights[50][48] = 16'sd-55;
        fc2_weights[50][49] = 16'sd-62;
        fc2_weights[50][50] = 16'sd6;
        fc2_weights[50][51] = 16'sd-33;
        fc2_weights[50][52] = 16'sd-17;
        fc2_weights[50][53] = 16'sd-20;
        fc2_weights[50][54] = 16'sd-69;
        fc2_weights[50][55] = 16'sd-15;
        fc2_weights[50][56] = 16'sd-26;
        fc2_weights[50][57] = 16'sd-43;
        fc2_weights[50][58] = 16'sd-5;
        fc2_weights[50][59] = 16'sd52;
        fc2_weights[50][60] = 16'sd-10;
        fc2_weights[50][61] = 16'sd51;
        fc2_weights[50][62] = 16'sd-100;
        fc2_weights[50][63] = 16'sd7;
        fc2_weights[50][64] = 16'sd-42;
        fc2_weights[50][65] = 16'sd-37;
        fc2_weights[50][66] = 16'sd-98;
        fc2_weights[50][67] = 16'sd9;
        fc2_weights[50][68] = 16'sd83;
        fc2_weights[50][69] = 16'sd-19;
        fc2_weights[50][70] = 16'sd-55;
        fc2_weights[50][71] = 16'sd-32;
        fc2_weights[50][72] = 16'sd-2;
        fc2_weights[50][73] = 16'sd10;
        fc2_weights[50][74] = 16'sd-27;
        fc2_weights[50][75] = 16'sd32;
        fc2_weights[50][76] = 16'sd-68;
        fc2_weights[50][77] = 16'sd-41;
        fc2_weights[50][78] = 16'sd-15;
        fc2_weights[50][79] = 16'sd29;
        fc2_weights[50][80] = 16'sd1;
        fc2_weights[50][81] = 16'sd-99;
        fc2_weights[50][82] = 16'sd7;
        fc2_weights[50][83] = 16'sd-30;
        fc2_weights[50][84] = 16'sd-20;
        fc2_weights[50][85] = 16'sd-3;
        fc2_weights[50][86] = 16'sd-71;
        fc2_weights[50][87] = 16'sd36;
        fc2_weights[50][88] = 16'sd7;
        fc2_weights[50][89] = 16'sd23;
        fc2_weights[50][90] = 16'sd-17;
        fc2_weights[50][91] = 16'sd-67;
        fc2_weights[50][92] = 16'sd-39;
        fc2_weights[50][93] = 16'sd26;
        fc2_weights[50][94] = 16'sd8;
        fc2_weights[50][95] = 16'sd-54;
        fc2_weights[50][96] = 16'sd-38;
        fc2_weights[50][97] = 16'sd15;
        fc2_weights[50][98] = 16'sd-9;
        fc2_weights[50][99] = 16'sd47;
        fc2_weights[50][100] = 16'sd-8;
        fc2_weights[50][101] = 16'sd6;
        fc2_weights[50][102] = 16'sd-77;
        fc2_weights[50][103] = 16'sd-15;
        fc2_weights[50][104] = 16'sd-12;
        fc2_weights[50][105] = 16'sd-11;
        fc2_weights[50][106] = 16'sd15;
        fc2_weights[50][107] = 16'sd-30;
        fc2_weights[50][108] = 16'sd-68;
        fc2_weights[50][109] = 16'sd-5;
        fc2_weights[50][110] = 16'sd-3;
        fc2_weights[50][111] = 16'sd7;
        fc2_weights[50][112] = 16'sd26;
        fc2_weights[50][113] = 16'sd31;
        fc2_weights[50][114] = 16'sd-69;
        fc2_weights[50][115] = 16'sd-15;
        fc2_weights[50][116] = 16'sd1;
        fc2_weights[50][117] = 16'sd-36;
        fc2_weights[50][118] = 16'sd9;
        fc2_weights[50][119] = 16'sd-30;
        fc2_weights[50][120] = 16'sd84;
        fc2_weights[50][121] = 16'sd-4;
        fc2_weights[50][122] = 16'sd-8;
        fc2_weights[50][123] = 16'sd-43;
        fc2_weights[50][124] = 16'sd80;
        fc2_weights[50][125] = 16'sd-29;
        fc2_weights[50][126] = 16'sd-52;
        fc2_weights[50][127] = 16'sd1;
        fc2_weights[51][0] = 16'sd39;
        fc2_weights[51][1] = 16'sd-19;
        fc2_weights[51][2] = 16'sd-11;
        fc2_weights[51][3] = 16'sd66;
        fc2_weights[51][4] = 16'sd22;
        fc2_weights[51][5] = 16'sd-10;
        fc2_weights[51][6] = 16'sd25;
        fc2_weights[51][7] = 16'sd-9;
        fc2_weights[51][8] = 16'sd32;
        fc2_weights[51][9] = 16'sd27;
        fc2_weights[51][10] = 16'sd-27;
        fc2_weights[51][11] = 16'sd-18;
        fc2_weights[51][12] = 16'sd66;
        fc2_weights[51][13] = 16'sd-34;
        fc2_weights[51][14] = 16'sd-81;
        fc2_weights[51][15] = 16'sd11;
        fc2_weights[51][16] = 16'sd2;
        fc2_weights[51][17] = 16'sd12;
        fc2_weights[51][18] = 16'sd-7;
        fc2_weights[51][19] = 16'sd-37;
        fc2_weights[51][20] = 16'sd14;
        fc2_weights[51][21] = 16'sd0;
        fc2_weights[51][22] = 16'sd-11;
        fc2_weights[51][23] = 16'sd15;
        fc2_weights[51][24] = 16'sd-24;
        fc2_weights[51][25] = 16'sd-24;
        fc2_weights[51][26] = 16'sd11;
        fc2_weights[51][27] = 16'sd-17;
        fc2_weights[51][28] = 16'sd21;
        fc2_weights[51][29] = 16'sd-20;
        fc2_weights[51][30] = 16'sd33;
        fc2_weights[51][31] = 16'sd21;
        fc2_weights[51][32] = 16'sd47;
        fc2_weights[51][33] = 16'sd41;
        fc2_weights[51][34] = 16'sd-32;
        fc2_weights[51][35] = 16'sd-66;
        fc2_weights[51][36] = 16'sd13;
        fc2_weights[51][37] = 16'sd-15;
        fc2_weights[51][38] = 16'sd74;
        fc2_weights[51][39] = 16'sd47;
        fc2_weights[51][40] = 16'sd-11;
        fc2_weights[51][41] = 16'sd-34;
        fc2_weights[51][42] = 16'sd-13;
        fc2_weights[51][43] = 16'sd28;
        fc2_weights[51][44] = 16'sd-45;
        fc2_weights[51][45] = 16'sd-88;
        fc2_weights[51][46] = 16'sd-46;
        fc2_weights[51][47] = 16'sd-6;
        fc2_weights[51][48] = 16'sd-27;
        fc2_weights[51][49] = 16'sd-22;
        fc2_weights[51][50] = 16'sd-55;
        fc2_weights[51][51] = 16'sd-41;
        fc2_weights[51][52] = 16'sd-65;
        fc2_weights[51][53] = 16'sd74;
        fc2_weights[51][54] = 16'sd-71;
        fc2_weights[51][55] = 16'sd-9;
        fc2_weights[51][56] = 16'sd-40;
        fc2_weights[51][57] = 16'sd-45;
        fc2_weights[51][58] = 16'sd-53;
        fc2_weights[51][59] = 16'sd16;
        fc2_weights[51][60] = 16'sd-75;
        fc2_weights[51][61] = 16'sd8;
        fc2_weights[51][62] = 16'sd-68;
        fc2_weights[51][63] = 16'sd-30;
        fc2_weights[51][64] = 16'sd11;
        fc2_weights[51][65] = 16'sd-47;
        fc2_weights[51][66] = 16'sd-27;
        fc2_weights[51][67] = 16'sd-7;
        fc2_weights[51][68] = 16'sd59;
        fc2_weights[51][69] = 16'sd-20;
        fc2_weights[51][70] = 16'sd24;
        fc2_weights[51][71] = 16'sd-43;
        fc2_weights[51][72] = 16'sd18;
        fc2_weights[51][73] = 16'sd6;
        fc2_weights[51][74] = 16'sd-52;
        fc2_weights[51][75] = 16'sd-29;
        fc2_weights[51][76] = 16'sd-37;
        fc2_weights[51][77] = 16'sd-61;
        fc2_weights[51][78] = 16'sd-18;
        fc2_weights[51][79] = 16'sd30;
        fc2_weights[51][80] = 16'sd47;
        fc2_weights[51][81] = 16'sd-55;
        fc2_weights[51][82] = 16'sd13;
        fc2_weights[51][83] = 16'sd-18;
        fc2_weights[51][84] = 16'sd35;
        fc2_weights[51][85] = 16'sd11;
        fc2_weights[51][86] = 16'sd23;
        fc2_weights[51][87] = 16'sd-8;
        fc2_weights[51][88] = 16'sd-12;
        fc2_weights[51][89] = 16'sd1;
        fc2_weights[51][90] = 16'sd-43;
        fc2_weights[51][91] = 16'sd-34;
        fc2_weights[51][92] = 16'sd-42;
        fc2_weights[51][93] = 16'sd68;
        fc2_weights[51][94] = 16'sd-11;
        fc2_weights[51][95] = 16'sd-11;
        fc2_weights[51][96] = 16'sd-5;
        fc2_weights[51][97] = 16'sd-35;
        fc2_weights[51][98] = 16'sd10;
        fc2_weights[51][99] = 16'sd17;
        fc2_weights[51][100] = 16'sd-74;
        fc2_weights[51][101] = 16'sd48;
        fc2_weights[51][102] = 16'sd-58;
        fc2_weights[51][103] = 16'sd-67;
        fc2_weights[51][104] = 16'sd-97;
        fc2_weights[51][105] = 16'sd-15;
        fc2_weights[51][106] = 16'sd36;
        fc2_weights[51][107] = 16'sd-19;
        fc2_weights[51][108] = 16'sd53;
        fc2_weights[51][109] = 16'sd48;
        fc2_weights[51][110] = 16'sd-31;
        fc2_weights[51][111] = 16'sd7;
        fc2_weights[51][112] = 16'sd17;
        fc2_weights[51][113] = 16'sd26;
        fc2_weights[51][114] = 16'sd-41;
        fc2_weights[51][115] = 16'sd20;
        fc2_weights[51][116] = 16'sd14;
        fc2_weights[51][117] = 16'sd8;
        fc2_weights[51][118] = 16'sd57;
        fc2_weights[51][119] = 16'sd-31;
        fc2_weights[51][120] = 16'sd48;
        fc2_weights[51][121] = 16'sd-24;
        fc2_weights[51][122] = 16'sd-79;
        fc2_weights[51][123] = 16'sd-81;
        fc2_weights[51][124] = 16'sd42;
        fc2_weights[51][125] = 16'sd-48;
        fc2_weights[51][126] = 16'sd-60;
        fc2_weights[51][127] = 16'sd-28;
        fc2_weights[52][0] = 16'sd-37;
        fc2_weights[52][1] = 16'sd-59;
        fc2_weights[52][2] = 16'sd61;
        fc2_weights[52][3] = 16'sd16;
        fc2_weights[52][4] = 16'sd-63;
        fc2_weights[52][5] = 16'sd-6;
        fc2_weights[52][6] = 16'sd-42;
        fc2_weights[52][7] = 16'sd-14;
        fc2_weights[52][8] = 16'sd-74;
        fc2_weights[52][9] = 16'sd-4;
        fc2_weights[52][10] = 16'sd-21;
        fc2_weights[52][11] = 16'sd-52;
        fc2_weights[52][12] = 16'sd-8;
        fc2_weights[52][13] = 16'sd34;
        fc2_weights[52][14] = 16'sd6;
        fc2_weights[52][15] = 16'sd18;
        fc2_weights[52][16] = 16'sd-1;
        fc2_weights[52][17] = 16'sd8;
        fc2_weights[52][18] = 16'sd-41;
        fc2_weights[52][19] = 16'sd42;
        fc2_weights[52][20] = 16'sd7;
        fc2_weights[52][21] = 16'sd-27;
        fc2_weights[52][22] = 16'sd-15;
        fc2_weights[52][23] = 16'sd-50;
        fc2_weights[52][24] = 16'sd18;
        fc2_weights[52][25] = 16'sd-16;
        fc2_weights[52][26] = 16'sd-2;
        fc2_weights[52][27] = 16'sd5;
        fc2_weights[52][28] = 16'sd-12;
        fc2_weights[52][29] = 16'sd-51;
        fc2_weights[52][30] = 16'sd20;
        fc2_weights[52][31] = 16'sd-20;
        fc2_weights[52][32] = 16'sd-17;
        fc2_weights[52][33] = 16'sd-20;
        fc2_weights[52][34] = 16'sd43;
        fc2_weights[52][35] = 16'sd37;
        fc2_weights[52][36] = 16'sd-67;
        fc2_weights[52][37] = 16'sd-5;
        fc2_weights[52][38] = 16'sd-14;
        fc2_weights[52][39] = 16'sd-9;
        fc2_weights[52][40] = 16'sd25;
        fc2_weights[52][41] = 16'sd35;
        fc2_weights[52][42] = 16'sd-7;
        fc2_weights[52][43] = 16'sd-28;
        fc2_weights[52][44] = 16'sd17;
        fc2_weights[52][45] = 16'sd87;
        fc2_weights[52][46] = 16'sd38;
        fc2_weights[52][47] = 16'sd-41;
        fc2_weights[52][48] = 16'sd40;
        fc2_weights[52][49] = 16'sd-26;
        fc2_weights[52][50] = 16'sd31;
        fc2_weights[52][51] = 16'sd-21;
        fc2_weights[52][52] = 16'sd20;
        fc2_weights[52][53] = 16'sd-85;
        fc2_weights[52][54] = 16'sd-53;
        fc2_weights[52][55] = 16'sd-7;
        fc2_weights[52][56] = 16'sd12;
        fc2_weights[52][57] = 16'sd25;
        fc2_weights[52][58] = 16'sd22;
        fc2_weights[52][59] = 16'sd-4;
        fc2_weights[52][60] = 16'sd-19;
        fc2_weights[52][61] = 16'sd-36;
        fc2_weights[52][62] = 16'sd8;
        fc2_weights[52][63] = 16'sd15;
        fc2_weights[52][64] = 16'sd-48;
        fc2_weights[52][65] = 16'sd0;
        fc2_weights[52][66] = 16'sd43;
        fc2_weights[52][67] = 16'sd-35;
        fc2_weights[52][68] = 16'sd-1;
        fc2_weights[52][69] = 16'sd11;
        fc2_weights[52][70] = 16'sd-32;
        fc2_weights[52][71] = 16'sd36;
        fc2_weights[52][72] = 16'sd-15;
        fc2_weights[52][73] = 16'sd-49;
        fc2_weights[52][74] = 16'sd-5;
        fc2_weights[52][75] = 16'sd-12;
        fc2_weights[52][76] = 16'sd19;
        fc2_weights[52][77] = 16'sd37;
        fc2_weights[52][78] = 16'sd15;
        fc2_weights[52][79] = 16'sd-18;
        fc2_weights[52][80] = 16'sd-78;
        fc2_weights[52][81] = 16'sd-24;
        fc2_weights[52][82] = 16'sd-39;
        fc2_weights[52][83] = 16'sd-16;
        fc2_weights[52][84] = 16'sd9;
        fc2_weights[52][85] = 16'sd-33;
        fc2_weights[52][86] = 16'sd-26;
        fc2_weights[52][87] = 16'sd-44;
        fc2_weights[52][88] = 16'sd22;
        fc2_weights[52][89] = 16'sd-83;
        fc2_weights[52][90] = 16'sd29;
        fc2_weights[52][91] = 16'sd-21;
        fc2_weights[52][92] = 16'sd-15;
        fc2_weights[52][93] = 16'sd-33;
        fc2_weights[52][94] = 16'sd43;
        fc2_weights[52][95] = 16'sd-50;
        fc2_weights[52][96] = 16'sd55;
        fc2_weights[52][97] = 16'sd-14;
        fc2_weights[52][98] = 16'sd-31;
        fc2_weights[52][99] = 16'sd-43;
        fc2_weights[52][100] = 16'sd24;
        fc2_weights[52][101] = 16'sd-24;
        fc2_weights[52][102] = 16'sd37;
        fc2_weights[52][103] = 16'sd50;
        fc2_weights[52][104] = 16'sd77;
        fc2_weights[52][105] = 16'sd-33;
        fc2_weights[52][106] = 16'sd-17;
        fc2_weights[52][107] = 16'sd13;
        fc2_weights[52][108] = 16'sd-68;
        fc2_weights[52][109] = 16'sd23;
        fc2_weights[52][110] = 16'sd-1;
        fc2_weights[52][111] = 16'sd-13;
        fc2_weights[52][112] = 16'sd-38;
        fc2_weights[52][113] = 16'sd-78;
        fc2_weights[52][114] = 16'sd-57;
        fc2_weights[52][115] = 16'sd-30;
        fc2_weights[52][116] = 16'sd55;
        fc2_weights[52][117] = 16'sd23;
        fc2_weights[52][118] = 16'sd-51;
        fc2_weights[52][119] = 16'sd-6;
        fc2_weights[52][120] = 16'sd-46;
        fc2_weights[52][121] = 16'sd-9;
        fc2_weights[52][122] = 16'sd0;
        fc2_weights[52][123] = 16'sd32;
        fc2_weights[52][124] = 16'sd-46;
        fc2_weights[52][125] = 16'sd71;
        fc2_weights[52][126] = 16'sd15;
        fc2_weights[52][127] = 16'sd31;
        fc2_weights[53][0] = 16'sd28;
        fc2_weights[53][1] = 16'sd-55;
        fc2_weights[53][2] = 16'sd-31;
        fc2_weights[53][3] = 16'sd-2;
        fc2_weights[53][4] = 16'sd30;
        fc2_weights[53][5] = 16'sd63;
        fc2_weights[53][6] = 16'sd-15;
        fc2_weights[53][7] = 16'sd-16;
        fc2_weights[53][8] = 16'sd-40;
        fc2_weights[53][9] = 16'sd-2;
        fc2_weights[53][10] = 16'sd23;
        fc2_weights[53][11] = 16'sd12;
        fc2_weights[53][12] = 16'sd-32;
        fc2_weights[53][13] = 16'sd16;
        fc2_weights[53][14] = 16'sd3;
        fc2_weights[53][15] = 16'sd-28;
        fc2_weights[53][16] = 16'sd87;
        fc2_weights[53][17] = 16'sd-44;
        fc2_weights[53][18] = 16'sd-37;
        fc2_weights[53][19] = 16'sd-77;
        fc2_weights[53][20] = 16'sd-76;
        fc2_weights[53][21] = 16'sd53;
        fc2_weights[53][22] = 16'sd-74;
        fc2_weights[53][23] = 16'sd22;
        fc2_weights[53][24] = 16'sd-63;
        fc2_weights[53][25] = 16'sd47;
        fc2_weights[53][26] = 16'sd6;
        fc2_weights[53][27] = 16'sd9;
        fc2_weights[53][28] = 16'sd33;
        fc2_weights[53][29] = 16'sd-17;
        fc2_weights[53][30] = 16'sd3;
        fc2_weights[53][31] = 16'sd33;
        fc2_weights[53][32] = 16'sd-48;
        fc2_weights[53][33] = 16'sd-19;
        fc2_weights[53][34] = 16'sd-73;
        fc2_weights[53][35] = 16'sd59;
        fc2_weights[53][36] = 16'sd-61;
        fc2_weights[53][37] = 16'sd-47;
        fc2_weights[53][38] = 16'sd3;
        fc2_weights[53][39] = 16'sd-3;
        fc2_weights[53][40] = 16'sd12;
        fc2_weights[53][41] = 16'sd-41;
        fc2_weights[53][42] = 16'sd-5;
        fc2_weights[53][43] = 16'sd-36;
        fc2_weights[53][44] = 16'sd-1;
        fc2_weights[53][45] = 16'sd59;
        fc2_weights[53][46] = 16'sd19;
        fc2_weights[53][47] = 16'sd-57;
        fc2_weights[53][48] = 16'sd20;
        fc2_weights[53][49] = 16'sd-29;
        fc2_weights[53][50] = 16'sd-5;
        fc2_weights[53][51] = 16'sd7;
        fc2_weights[53][52] = 16'sd-103;
        fc2_weights[53][53] = 16'sd-30;
        fc2_weights[53][54] = 16'sd10;
        fc2_weights[53][55] = 16'sd46;
        fc2_weights[53][56] = 16'sd29;
        fc2_weights[53][57] = 16'sd-34;
        fc2_weights[53][58] = 16'sd-29;
        fc2_weights[53][59] = 16'sd-67;
        fc2_weights[53][60] = 16'sd-59;
        fc2_weights[53][61] = 16'sd23;
        fc2_weights[53][62] = 16'sd-51;
        fc2_weights[53][63] = 16'sd-37;
        fc2_weights[53][64] = 16'sd-44;
        fc2_weights[53][65] = 16'sd-78;
        fc2_weights[53][66] = 16'sd3;
        fc2_weights[53][67] = 16'sd13;
        fc2_weights[53][68] = 16'sd-76;
        fc2_weights[53][69] = 16'sd18;
        fc2_weights[53][70] = 16'sd27;
        fc2_weights[53][71] = 16'sd1;
        fc2_weights[53][72] = 16'sd52;
        fc2_weights[53][73] = 16'sd-19;
        fc2_weights[53][74] = 16'sd-31;
        fc2_weights[53][75] = 16'sd59;
        fc2_weights[53][76] = 16'sd37;
        fc2_weights[53][77] = 16'sd-35;
        fc2_weights[53][78] = 16'sd16;
        fc2_weights[53][79] = 16'sd-5;
        fc2_weights[53][80] = 16'sd-21;
        fc2_weights[53][81] = 16'sd-15;
        fc2_weights[53][82] = 16'sd0;
        fc2_weights[53][83] = 16'sd54;
        fc2_weights[53][84] = 16'sd-72;
        fc2_weights[53][85] = 16'sd9;
        fc2_weights[53][86] = 16'sd-14;
        fc2_weights[53][87] = 16'sd-50;
        fc2_weights[53][88] = 16'sd23;
        fc2_weights[53][89] = 16'sd45;
        fc2_weights[53][90] = 16'sd-22;
        fc2_weights[53][91] = 16'sd53;
        fc2_weights[53][92] = 16'sd-28;
        fc2_weights[53][93] = 16'sd-54;
        fc2_weights[53][94] = 16'sd-66;
        fc2_weights[53][95] = 16'sd32;
        fc2_weights[53][96] = 16'sd-11;
        fc2_weights[53][97] = 16'sd-55;
        fc2_weights[53][98] = 16'sd71;
        fc2_weights[53][99] = 16'sd-65;
        fc2_weights[53][100] = 16'sd-42;
        fc2_weights[53][101] = 16'sd-27;
        fc2_weights[53][102] = 16'sd19;
        fc2_weights[53][103] = 16'sd6;
        fc2_weights[53][104] = 16'sd-36;
        fc2_weights[53][105] = 16'sd-13;
        fc2_weights[53][106] = 16'sd18;
        fc2_weights[53][107] = 16'sd27;
        fc2_weights[53][108] = 16'sd-53;
        fc2_weights[53][109] = 16'sd-38;
        fc2_weights[53][110] = 16'sd42;
        fc2_weights[53][111] = 16'sd-14;
        fc2_weights[53][112] = 16'sd0;
        fc2_weights[53][113] = 16'sd-16;
        fc2_weights[53][114] = 16'sd48;
        fc2_weights[53][115] = 16'sd26;
        fc2_weights[53][116] = 16'sd2;
        fc2_weights[53][117] = 16'sd-74;
        fc2_weights[53][118] = 16'sd-26;
        fc2_weights[53][119] = 16'sd-6;
        fc2_weights[53][120] = 16'sd-38;
        fc2_weights[53][121] = 16'sd-11;
        fc2_weights[53][122] = 16'sd40;
        fc2_weights[53][123] = 16'sd23;
        fc2_weights[53][124] = 16'sd-44;
        fc2_weights[53][125] = 16'sd-16;
        fc2_weights[53][126] = 16'sd-40;
        fc2_weights[53][127] = 16'sd-8;
        fc2_weights[54][0] = 16'sd17;
        fc2_weights[54][1] = 16'sd3;
        fc2_weights[54][2] = 16'sd-14;
        fc2_weights[54][3] = 16'sd-14;
        fc2_weights[54][4] = 16'sd-40;
        fc2_weights[54][5] = 16'sd52;
        fc2_weights[54][6] = 16'sd60;
        fc2_weights[54][7] = 16'sd23;
        fc2_weights[54][8] = 16'sd52;
        fc2_weights[54][9] = 16'sd29;
        fc2_weights[54][10] = 16'sd-11;
        fc2_weights[54][11] = 16'sd7;
        fc2_weights[54][12] = 16'sd86;
        fc2_weights[54][13] = 16'sd-43;
        fc2_weights[54][14] = 16'sd-25;
        fc2_weights[54][15] = 16'sd12;
        fc2_weights[54][16] = 16'sd-37;
        fc2_weights[54][17] = 16'sd26;
        fc2_weights[54][18] = 16'sd25;
        fc2_weights[54][19] = 16'sd22;
        fc2_weights[54][20] = 16'sd32;
        fc2_weights[54][21] = 16'sd3;
        fc2_weights[54][22] = 16'sd-7;
        fc2_weights[54][23] = 16'sd-5;
        fc2_weights[54][24] = 16'sd-32;
        fc2_weights[54][25] = 16'sd-20;
        fc2_weights[54][26] = 16'sd-6;
        fc2_weights[54][27] = 16'sd-19;
        fc2_weights[54][28] = 16'sd65;
        fc2_weights[54][29] = 16'sd-24;
        fc2_weights[54][30] = 16'sd22;
        fc2_weights[54][31] = 16'sd33;
        fc2_weights[54][32] = 16'sd-1;
        fc2_weights[54][33] = 16'sd83;
        fc2_weights[54][34] = 16'sd-6;
        fc2_weights[54][35] = 16'sd-56;
        fc2_weights[54][36] = 16'sd24;
        fc2_weights[54][37] = 16'sd23;
        fc2_weights[54][38] = 16'sd-43;
        fc2_weights[54][39] = 16'sd59;
        fc2_weights[54][40] = 16'sd-55;
        fc2_weights[54][41] = 16'sd-60;
        fc2_weights[54][42] = 16'sd-65;
        fc2_weights[54][43] = 16'sd59;
        fc2_weights[54][44] = 16'sd-8;
        fc2_weights[54][45] = 16'sd-73;
        fc2_weights[54][46] = 16'sd-39;
        fc2_weights[54][47] = 16'sd34;
        fc2_weights[54][48] = 16'sd-54;
        fc2_weights[54][49] = 16'sd-58;
        fc2_weights[54][50] = 16'sd-46;
        fc2_weights[54][51] = 16'sd-107;
        fc2_weights[54][52] = 16'sd-16;
        fc2_weights[54][53] = 16'sd87;
        fc2_weights[54][54] = 16'sd-19;
        fc2_weights[54][55] = 16'sd44;
        fc2_weights[54][56] = 16'sd-21;
        fc2_weights[54][57] = 16'sd-62;
        fc2_weights[54][58] = 16'sd25;
        fc2_weights[54][59] = 16'sd25;
        fc2_weights[54][60] = 16'sd-67;
        fc2_weights[54][61] = 16'sd2;
        fc2_weights[54][62] = 16'sd-45;
        fc2_weights[54][63] = 16'sd-9;
        fc2_weights[54][64] = 16'sd44;
        fc2_weights[54][65] = 16'sd-45;
        fc2_weights[54][66] = 16'sd-50;
        fc2_weights[54][67] = 16'sd-14;
        fc2_weights[54][68] = 16'sd111;
        fc2_weights[54][69] = 16'sd7;
        fc2_weights[54][70] = 16'sd-10;
        fc2_weights[54][71] = 16'sd-47;
        fc2_weights[54][72] = 16'sd59;
        fc2_weights[54][73] = 16'sd19;
        fc2_weights[54][74] = 16'sd-12;
        fc2_weights[54][75] = 16'sd-43;
        fc2_weights[54][76] = 16'sd-36;
        fc2_weights[54][77] = 16'sd-71;
        fc2_weights[54][78] = 16'sd-28;
        fc2_weights[54][79] = 16'sd-5;
        fc2_weights[54][80] = 16'sd63;
        fc2_weights[54][81] = 16'sd-32;
        fc2_weights[54][82] = 16'sd35;
        fc2_weights[54][83] = 16'sd-58;
        fc2_weights[54][84] = 16'sd-16;
        fc2_weights[54][85] = 16'sd-26;
        fc2_weights[54][86] = 16'sd-39;
        fc2_weights[54][87] = 16'sd41;
        fc2_weights[54][88] = 16'sd4;
        fc2_weights[54][89] = 16'sd37;
        fc2_weights[54][90] = 16'sd-47;
        fc2_weights[54][91] = 16'sd-12;
        fc2_weights[54][92] = 16'sd-49;
        fc2_weights[54][93] = 16'sd46;
        fc2_weights[54][94] = 16'sd17;
        fc2_weights[54][95] = 16'sd20;
        fc2_weights[54][96] = 16'sd-44;
        fc2_weights[54][97] = 16'sd-36;
        fc2_weights[54][98] = 16'sd-66;
        fc2_weights[54][99] = 16'sd10;
        fc2_weights[54][100] = 16'sd-101;
        fc2_weights[54][101] = 16'sd76;
        fc2_weights[54][102] = 16'sd-45;
        fc2_weights[54][103] = 16'sd-73;
        fc2_weights[54][104] = 16'sd-69;
        fc2_weights[54][105] = 16'sd-15;
        fc2_weights[54][106] = 16'sd0;
        fc2_weights[54][107] = 16'sd-28;
        fc2_weights[54][108] = 16'sd41;
        fc2_weights[54][109] = 16'sd-14;
        fc2_weights[54][110] = 16'sd-42;
        fc2_weights[54][111] = 16'sd-17;
        fc2_weights[54][112] = 16'sd35;
        fc2_weights[54][113] = 16'sd51;
        fc2_weights[54][114] = 16'sd-22;
        fc2_weights[54][115] = 16'sd1;
        fc2_weights[54][116] = 16'sd-1;
        fc2_weights[54][117] = 16'sd-25;
        fc2_weights[54][118] = 16'sd24;
        fc2_weights[54][119] = 16'sd8;
        fc2_weights[54][120] = 16'sd58;
        fc2_weights[54][121] = 16'sd1;
        fc2_weights[54][122] = 16'sd-52;
        fc2_weights[54][123] = 16'sd-44;
        fc2_weights[54][124] = 16'sd37;
        fc2_weights[54][125] = 16'sd-20;
        fc2_weights[54][126] = 16'sd-94;
        fc2_weights[54][127] = 16'sd-52;
        fc2_weights[55][0] = 16'sd54;
        fc2_weights[55][1] = 16'sd-2;
        fc2_weights[55][2] = 16'sd-10;
        fc2_weights[55][3] = 16'sd71;
        fc2_weights[55][4] = 16'sd10;
        fc2_weights[55][5] = 16'sd5;
        fc2_weights[55][6] = 16'sd6;
        fc2_weights[55][7] = 16'sd-13;
        fc2_weights[55][8] = 16'sd15;
        fc2_weights[55][9] = 16'sd30;
        fc2_weights[55][10] = 16'sd-20;
        fc2_weights[55][11] = 16'sd-16;
        fc2_weights[55][12] = 16'sd6;
        fc2_weights[55][13] = 16'sd43;
        fc2_weights[55][14] = 16'sd-30;
        fc2_weights[55][15] = 16'sd2;
        fc2_weights[55][16] = 16'sd1;
        fc2_weights[55][17] = 16'sd78;
        fc2_weights[55][18] = 16'sd-2;
        fc2_weights[55][19] = 16'sd-3;
        fc2_weights[55][20] = 16'sd19;
        fc2_weights[55][21] = 16'sd-32;
        fc2_weights[55][22] = 16'sd-39;
        fc2_weights[55][23] = 16'sd-42;
        fc2_weights[55][24] = 16'sd-2;
        fc2_weights[55][25] = 16'sd-31;
        fc2_weights[55][26] = 16'sd-8;
        fc2_weights[55][27] = 16'sd6;
        fc2_weights[55][28] = 16'sd-21;
        fc2_weights[55][29] = 16'sd-30;
        fc2_weights[55][30] = 16'sd33;
        fc2_weights[55][31] = 16'sd-27;
        fc2_weights[55][32] = 16'sd-12;
        fc2_weights[55][33] = 16'sd13;
        fc2_weights[55][34] = 16'sd22;
        fc2_weights[55][35] = 16'sd15;
        fc2_weights[55][36] = 16'sd-25;
        fc2_weights[55][37] = 16'sd-34;
        fc2_weights[55][38] = 16'sd1;
        fc2_weights[55][39] = 16'sd-7;
        fc2_weights[55][40] = 16'sd15;
        fc2_weights[55][41] = 16'sd-7;
        fc2_weights[55][42] = 16'sd32;
        fc2_weights[55][43] = 16'sd-16;
        fc2_weights[55][44] = 16'sd37;
        fc2_weights[55][45] = 16'sd27;
        fc2_weights[55][46] = 16'sd-42;
        fc2_weights[55][47] = 16'sd-35;
        fc2_weights[55][48] = 16'sd73;
        fc2_weights[55][49] = 16'sd-11;
        fc2_weights[55][50] = 16'sd79;
        fc2_weights[55][51] = 16'sd-5;
        fc2_weights[55][52] = 16'sd51;
        fc2_weights[55][53] = 16'sd-23;
        fc2_weights[55][54] = 16'sd-52;
        fc2_weights[55][55] = 16'sd4;
        fc2_weights[55][56] = 16'sd26;
        fc2_weights[55][57] = 16'sd-20;
        fc2_weights[55][58] = 16'sd24;
        fc2_weights[55][59] = 16'sd4;
        fc2_weights[55][60] = 16'sd-25;
        fc2_weights[55][61] = 16'sd-11;
        fc2_weights[55][62] = 16'sd-2;
        fc2_weights[55][63] = 16'sd12;
        fc2_weights[55][64] = 16'sd-47;
        fc2_weights[55][65] = 16'sd58;
        fc2_weights[55][66] = 16'sd-39;
        fc2_weights[55][67] = 16'sd-24;
        fc2_weights[55][68] = 16'sd-7;
        fc2_weights[55][69] = 16'sd-5;
        fc2_weights[55][70] = 16'sd-54;
        fc2_weights[55][71] = 16'sd-18;
        fc2_weights[55][72] = 16'sd-6;
        fc2_weights[55][73] = 16'sd-14;
        fc2_weights[55][74] = 16'sd16;
        fc2_weights[55][75] = 16'sd3;
        fc2_weights[55][76] = 16'sd-61;
        fc2_weights[55][77] = 16'sd-19;
        fc2_weights[55][78] = 16'sd30;
        fc2_weights[55][79] = 16'sd-17;
        fc2_weights[55][80] = 16'sd-49;
        fc2_weights[55][81] = 16'sd2;
        fc2_weights[55][82] = 16'sd0;
        fc2_weights[55][83] = 16'sd-23;
        fc2_weights[55][84] = 16'sd-21;
        fc2_weights[55][85] = 16'sd36;
        fc2_weights[55][86] = 16'sd-10;
        fc2_weights[55][87] = 16'sd0;
        fc2_weights[55][88] = 16'sd21;
        fc2_weights[55][89] = 16'sd-5;
        fc2_weights[55][90] = 16'sd-1;
        fc2_weights[55][91] = 16'sd-30;
        fc2_weights[55][92] = 16'sd-30;
        fc2_weights[55][93] = 16'sd47;
        fc2_weights[55][94] = 16'sd10;
        fc2_weights[55][95] = 16'sd-31;
        fc2_weights[55][96] = 16'sd7;
        fc2_weights[55][97] = 16'sd12;
        fc2_weights[55][98] = 16'sd-40;
        fc2_weights[55][99] = 16'sd-7;
        fc2_weights[55][100] = 16'sd8;
        fc2_weights[55][101] = 16'sd-7;
        fc2_weights[55][102] = 16'sd-36;
        fc2_weights[55][103] = 16'sd52;
        fc2_weights[55][104] = 16'sd74;
        fc2_weights[55][105] = 16'sd6;
        fc2_weights[55][106] = 16'sd-24;
        fc2_weights[55][107] = 16'sd-24;
        fc2_weights[55][108] = 16'sd-12;
        fc2_weights[55][109] = 16'sd-34;
        fc2_weights[55][110] = 16'sd47;
        fc2_weights[55][111] = 16'sd-3;
        fc2_weights[55][112] = 16'sd-9;
        fc2_weights[55][113] = 16'sd-8;
        fc2_weights[55][114] = 16'sd-13;
        fc2_weights[55][115] = 16'sd-18;
        fc2_weights[55][116] = 16'sd3;
        fc2_weights[55][117] = 16'sd-2;
        fc2_weights[55][118] = 16'sd-31;
        fc2_weights[55][119] = 16'sd-20;
        fc2_weights[55][120] = 16'sd-39;
        fc2_weights[55][121] = 16'sd5;
        fc2_weights[55][122] = 16'sd3;
        fc2_weights[55][123] = 16'sd51;
        fc2_weights[55][124] = 16'sd6;
        fc2_weights[55][125] = 16'sd55;
        fc2_weights[55][126] = 16'sd17;
        fc2_weights[55][127] = 16'sd-10;
        fc2_weights[56][0] = 16'sd-48;
        fc2_weights[56][1] = 16'sd-22;
        fc2_weights[56][2] = 16'sd12;
        fc2_weights[56][3] = 16'sd-36;
        fc2_weights[56][4] = 16'sd-22;
        fc2_weights[56][5] = 16'sd24;
        fc2_weights[56][6] = 16'sd5;
        fc2_weights[56][7] = 16'sd-63;
        fc2_weights[56][8] = 16'sd54;
        fc2_weights[56][9] = 16'sd-10;
        fc2_weights[56][10] = 16'sd-18;
        fc2_weights[56][11] = 16'sd0;
        fc2_weights[56][12] = 16'sd11;
        fc2_weights[56][13] = 16'sd-7;
        fc2_weights[56][14] = 16'sd3;
        fc2_weights[56][15] = 16'sd-2;
        fc2_weights[56][16] = 16'sd23;
        fc2_weights[56][17] = 16'sd17;
        fc2_weights[56][18] = 16'sd-19;
        fc2_weights[56][19] = 16'sd-18;
        fc2_weights[56][20] = 16'sd17;
        fc2_weights[56][21] = 16'sd-45;
        fc2_weights[56][22] = 16'sd-79;
        fc2_weights[56][23] = 16'sd17;
        fc2_weights[56][24] = 16'sd-48;
        fc2_weights[56][25] = 16'sd31;
        fc2_weights[56][26] = 16'sd15;
        fc2_weights[56][27] = 16'sd6;
        fc2_weights[56][28] = 16'sd-25;
        fc2_weights[56][29] = 16'sd-4;
        fc2_weights[56][30] = 16'sd0;
        fc2_weights[56][31] = 16'sd7;
        fc2_weights[56][32] = 16'sd-9;
        fc2_weights[56][33] = 16'sd-3;
        fc2_weights[56][34] = 16'sd-9;
        fc2_weights[56][35] = 16'sd-49;
        fc2_weights[56][36] = 16'sd-37;
        fc2_weights[56][37] = 16'sd-1;
        fc2_weights[56][38] = 16'sd-16;
        fc2_weights[56][39] = 16'sd50;
        fc2_weights[56][40] = 16'sd-39;
        fc2_weights[56][41] = 16'sd113;
        fc2_weights[56][42] = 16'sd9;
        fc2_weights[56][43] = 16'sd-41;
        fc2_weights[56][44] = 16'sd7;
        fc2_weights[56][45] = 16'sd-18;
        fc2_weights[56][46] = 16'sd-50;
        fc2_weights[56][47] = 16'sd4;
        fc2_weights[56][48] = 16'sd34;
        fc2_weights[56][49] = 16'sd3;
        fc2_weights[56][50] = 16'sd8;
        fc2_weights[56][51] = 16'sd8;
        fc2_weights[56][52] = 16'sd-7;
        fc2_weights[56][53] = 16'sd20;
        fc2_weights[56][54] = 16'sd-1;
        fc2_weights[56][55] = 16'sd-7;
        fc2_weights[56][56] = 16'sd25;
        fc2_weights[56][57] = 16'sd-6;
        fc2_weights[56][58] = 16'sd23;
        fc2_weights[56][59] = 16'sd10;
        fc2_weights[56][60] = 16'sd15;
        fc2_weights[56][61] = 16'sd-35;
        fc2_weights[56][62] = 16'sd21;
        fc2_weights[56][63] = 16'sd-12;
        fc2_weights[56][64] = 16'sd-13;
        fc2_weights[56][65] = 16'sd10;
        fc2_weights[56][66] = 16'sd6;
        fc2_weights[56][67] = 16'sd-31;
        fc2_weights[56][68] = 16'sd-21;
        fc2_weights[56][69] = 16'sd12;
        fc2_weights[56][70] = 16'sd29;
        fc2_weights[56][71] = 16'sd30;
        fc2_weights[56][72] = 16'sd68;
        fc2_weights[56][73] = 16'sd-20;
        fc2_weights[56][74] = 16'sd-32;
        fc2_weights[56][75] = 16'sd28;
        fc2_weights[56][76] = 16'sd8;
        fc2_weights[56][77] = 16'sd36;
        fc2_weights[56][78] = 16'sd33;
        fc2_weights[56][79] = 16'sd-6;
        fc2_weights[56][80] = 16'sd15;
        fc2_weights[56][81] = 16'sd-30;
        fc2_weights[56][82] = 16'sd-2;
        fc2_weights[56][83] = 16'sd23;
        fc2_weights[56][84] = 16'sd-1;
        fc2_weights[56][85] = 16'sd-11;
        fc2_weights[56][86] = 16'sd17;
        fc2_weights[56][87] = 16'sd-45;
        fc2_weights[56][88] = 16'sd20;
        fc2_weights[56][89] = 16'sd0;
        fc2_weights[56][90] = 16'sd-23;
        fc2_weights[56][91] = 16'sd24;
        fc2_weights[56][92] = 16'sd10;
        fc2_weights[56][93] = 16'sd-15;
        fc2_weights[56][94] = 16'sd-54;
        fc2_weights[56][95] = 16'sd14;
        fc2_weights[56][96] = 16'sd23;
        fc2_weights[56][97] = 16'sd132;
        fc2_weights[56][98] = 16'sd15;
        fc2_weights[56][99] = 16'sd12;
        fc2_weights[56][100] = 16'sd-20;
        fc2_weights[56][101] = 16'sd-27;
        fc2_weights[56][102] = 16'sd22;
        fc2_weights[56][103] = 16'sd-20;
        fc2_weights[56][104] = 16'sd2;
        fc2_weights[56][105] = 16'sd0;
        fc2_weights[56][106] = 16'sd-11;
        fc2_weights[56][107] = 16'sd70;
        fc2_weights[56][108] = 16'sd-28;
        fc2_weights[56][109] = 16'sd46;
        fc2_weights[56][110] = 16'sd34;
        fc2_weights[56][111] = 16'sd-4;
        fc2_weights[56][112] = 16'sd11;
        fc2_weights[56][113] = 16'sd12;
        fc2_weights[56][114] = 16'sd33;
        fc2_weights[56][115] = 16'sd46;
        fc2_weights[56][116] = 16'sd6;
        fc2_weights[56][117] = 16'sd-13;
        fc2_weights[56][118] = 16'sd8;
        fc2_weights[56][119] = 16'sd-11;
        fc2_weights[56][120] = 16'sd25;
        fc2_weights[56][121] = 16'sd86;
        fc2_weights[56][122] = 16'sd52;
        fc2_weights[56][123] = 16'sd-7;
        fc2_weights[56][124] = 16'sd32;
        fc2_weights[56][125] = 16'sd-24;
        fc2_weights[56][126] = 16'sd15;
        fc2_weights[56][127] = 16'sd-13;
        fc2_weights[57][0] = 16'sd42;
        fc2_weights[57][1] = 16'sd-30;
        fc2_weights[57][2] = 16'sd8;
        fc2_weights[57][3] = 16'sd-77;
        fc2_weights[57][4] = 16'sd24;
        fc2_weights[57][5] = 16'sd-29;
        fc2_weights[57][6] = 16'sd45;
        fc2_weights[57][7] = 16'sd-11;
        fc2_weights[57][8] = 16'sd11;
        fc2_weights[57][9] = 16'sd-31;
        fc2_weights[57][10] = 16'sd-5;
        fc2_weights[57][11] = 16'sd73;
        fc2_weights[57][12] = 16'sd-38;
        fc2_weights[57][13] = 16'sd-32;
        fc2_weights[57][14] = 16'sd41;
        fc2_weights[57][15] = 16'sd-37;
        fc2_weights[57][16] = 16'sd42;
        fc2_weights[57][17] = 16'sd-77;
        fc2_weights[57][18] = 16'sd-23;
        fc2_weights[57][19] = 16'sd-9;
        fc2_weights[57][20] = 16'sd-58;
        fc2_weights[57][21] = 16'sd-45;
        fc2_weights[57][22] = 16'sd15;
        fc2_weights[57][23] = 16'sd82;
        fc2_weights[57][24] = 16'sd-39;
        fc2_weights[57][25] = 16'sd-41;
        fc2_weights[57][26] = 16'sd35;
        fc2_weights[57][27] = 16'sd2;
        fc2_weights[57][28] = 16'sd11;
        fc2_weights[57][29] = 16'sd37;
        fc2_weights[57][30] = 16'sd-56;
        fc2_weights[57][31] = 16'sd22;
        fc2_weights[57][32] = 16'sd-52;
        fc2_weights[57][33] = 16'sd-32;
        fc2_weights[57][34] = 16'sd-23;
        fc2_weights[57][35] = 16'sd10;
        fc2_weights[57][36] = 16'sd16;
        fc2_weights[57][37] = 16'sd-53;
        fc2_weights[57][38] = 16'sd58;
        fc2_weights[57][39] = 16'sd-11;
        fc2_weights[57][40] = 16'sd-37;
        fc2_weights[57][41] = 16'sd41;
        fc2_weights[57][42] = 16'sd5;
        fc2_weights[57][43] = 16'sd-66;
        fc2_weights[57][44] = 16'sd33;
        fc2_weights[57][45] = 16'sd43;
        fc2_weights[57][46] = 16'sd72;
        fc2_weights[57][47] = 16'sd15;
        fc2_weights[57][48] = 16'sd-30;
        fc2_weights[57][49] = 16'sd29;
        fc2_weights[57][50] = 16'sd-22;
        fc2_weights[57][51] = 16'sd62;
        fc2_weights[57][52] = 16'sd-36;
        fc2_weights[57][53] = 16'sd17;
        fc2_weights[57][54] = 16'sd63;
        fc2_weights[57][55] = 16'sd-8;
        fc2_weights[57][56] = 16'sd17;
        fc2_weights[57][57] = 16'sd-58;
        fc2_weights[57][58] = 16'sd-34;
        fc2_weights[57][59] = 16'sd-35;
        fc2_weights[57][60] = 16'sd35;
        fc2_weights[57][61] = 16'sd-20;
        fc2_weights[57][62] = 16'sd62;
        fc2_weights[57][63] = 16'sd-18;
        fc2_weights[57][64] = 16'sd24;
        fc2_weights[57][65] = 16'sd-10;
        fc2_weights[57][66] = 16'sd8;
        fc2_weights[57][67] = 16'sd7;
        fc2_weights[57][68] = 16'sd-62;
        fc2_weights[57][69] = 16'sd-48;
        fc2_weights[57][70] = 16'sd54;
        fc2_weights[57][71] = 16'sd-11;
        fc2_weights[57][72] = 16'sd-7;
        fc2_weights[57][73] = 16'sd-22;
        fc2_weights[57][74] = 16'sd-16;
        fc2_weights[57][75] = 16'sd33;
        fc2_weights[57][76] = 16'sd-51;
        fc2_weights[57][77] = 16'sd89;
        fc2_weights[57][78] = 16'sd-64;
        fc2_weights[57][79] = 16'sd13;
        fc2_weights[57][80] = 16'sd8;
        fc2_weights[57][81] = 16'sd4;
        fc2_weights[57][82] = 16'sd-7;
        fc2_weights[57][83] = 16'sd37;
        fc2_weights[57][84] = 16'sd-17;
        fc2_weights[57][85] = 16'sd26;
        fc2_weights[57][86] = 16'sd4;
        fc2_weights[57][87] = 16'sd-37;
        fc2_weights[57][88] = 16'sd1;
        fc2_weights[57][89] = 16'sd18;
        fc2_weights[57][90] = 16'sd22;
        fc2_weights[57][91] = 16'sd8;
        fc2_weights[57][92] = 16'sd66;
        fc2_weights[57][93] = 16'sd18;
        fc2_weights[57][94] = 16'sd-80;
        fc2_weights[57][95] = 16'sd-3;
        fc2_weights[57][96] = 16'sd-30;
        fc2_weights[57][97] = 16'sd21;
        fc2_weights[57][98] = 16'sd50;
        fc2_weights[57][99] = 16'sd8;
        fc2_weights[57][100] = 16'sd5;
        fc2_weights[57][101] = 16'sd-64;
        fc2_weights[57][102] = 16'sd26;
        fc2_weights[57][103] = 16'sd-41;
        fc2_weights[57][104] = 16'sd59;
        fc2_weights[57][105] = 16'sd5;
        fc2_weights[57][106] = 16'sd11;
        fc2_weights[57][107] = 16'sd31;
        fc2_weights[57][108] = 16'sd-29;
        fc2_weights[57][109] = 16'sd11;
        fc2_weights[57][110] = 16'sd-3;
        fc2_weights[57][111] = 16'sd25;
        fc2_weights[57][112] = 16'sd-19;
        fc2_weights[57][113] = 16'sd-36;
        fc2_weights[57][114] = 16'sd0;
        fc2_weights[57][115] = 16'sd34;
        fc2_weights[57][116] = 16'sd25;
        fc2_weights[57][117] = 16'sd-81;
        fc2_weights[57][118] = 16'sd31;
        fc2_weights[57][119] = 16'sd-10;
        fc2_weights[57][120] = 16'sd-58;
        fc2_weights[57][121] = 16'sd3;
        fc2_weights[57][122] = 16'sd-17;
        fc2_weights[57][123] = 16'sd-6;
        fc2_weights[57][124] = 16'sd-42;
        fc2_weights[57][125] = 16'sd20;
        fc2_weights[57][126] = 16'sd29;
        fc2_weights[57][127] = 16'sd-47;
        fc2_weights[58][0] = 16'sd-57;
        fc2_weights[58][1] = 16'sd-49;
        fc2_weights[58][2] = 16'sd13;
        fc2_weights[58][3] = 16'sd34;
        fc2_weights[58][4] = 16'sd-91;
        fc2_weights[58][5] = 16'sd-23;
        fc2_weights[58][6] = 16'sd2;
        fc2_weights[58][7] = 16'sd24;
        fc2_weights[58][8] = 16'sd-69;
        fc2_weights[58][9] = 16'sd6;
        fc2_weights[58][10] = 16'sd17;
        fc2_weights[58][11] = 16'sd-35;
        fc2_weights[58][12] = 16'sd-24;
        fc2_weights[58][13] = 16'sd38;
        fc2_weights[58][14] = 16'sd4;
        fc2_weights[58][15] = 16'sd33;
        fc2_weights[58][16] = 16'sd22;
        fc2_weights[58][17] = 16'sd-8;
        fc2_weights[58][18] = 16'sd-53;
        fc2_weights[58][19] = 16'sd14;
        fc2_weights[58][20] = 16'sd20;
        fc2_weights[58][21] = 16'sd-23;
        fc2_weights[58][22] = 16'sd-48;
        fc2_weights[58][23] = 16'sd-47;
        fc2_weights[58][24] = 16'sd20;
        fc2_weights[58][25] = 16'sd-75;
        fc2_weights[58][26] = 16'sd46;
        fc2_weights[58][27] = 16'sd19;
        fc2_weights[58][28] = 16'sd-1;
        fc2_weights[58][29] = 16'sd-52;
        fc2_weights[58][30] = 16'sd-5;
        fc2_weights[58][31] = 16'sd-39;
        fc2_weights[58][32] = 16'sd30;
        fc2_weights[58][33] = 16'sd-5;
        fc2_weights[58][34] = 16'sd25;
        fc2_weights[58][35] = 16'sd44;
        fc2_weights[58][36] = 16'sd-57;
        fc2_weights[58][37] = 16'sd22;
        fc2_weights[58][38] = 16'sd-62;
        fc2_weights[58][39] = 16'sd-39;
        fc2_weights[58][40] = 16'sd37;
        fc2_weights[58][41] = 16'sd-18;
        fc2_weights[58][42] = 16'sd-25;
        fc2_weights[58][43] = 16'sd-23;
        fc2_weights[58][44] = 16'sd35;
        fc2_weights[58][45] = 16'sd3;
        fc2_weights[58][46] = 16'sd-14;
        fc2_weights[58][47] = 16'sd62;
        fc2_weights[58][48] = 16'sd-1;
        fc2_weights[58][49] = 16'sd-15;
        fc2_weights[58][50] = 16'sd19;
        fc2_weights[58][51] = 16'sd-10;
        fc2_weights[58][52] = 16'sd6;
        fc2_weights[58][53] = 16'sd-59;
        fc2_weights[58][54] = 16'sd11;
        fc2_weights[58][55] = 16'sd-55;
        fc2_weights[58][56] = 16'sd32;
        fc2_weights[58][57] = 16'sd67;
        fc2_weights[58][58] = 16'sd-1;
        fc2_weights[58][59] = 16'sd25;
        fc2_weights[58][60] = 16'sd16;
        fc2_weights[58][61] = 16'sd21;
        fc2_weights[58][62] = 16'sd-5;
        fc2_weights[58][63] = 16'sd46;
        fc2_weights[58][64] = 16'sd-5;
        fc2_weights[58][65] = 16'sd-11;
        fc2_weights[58][66] = 16'sd-16;
        fc2_weights[58][67] = 16'sd-51;
        fc2_weights[58][68] = 16'sd5;
        fc2_weights[58][69] = 16'sd66;
        fc2_weights[58][70] = 16'sd-27;
        fc2_weights[58][71] = 16'sd45;
        fc2_weights[58][72] = 16'sd-50;
        fc2_weights[58][73] = 16'sd-8;
        fc2_weights[58][74] = 16'sd20;
        fc2_weights[58][75] = 16'sd-3;
        fc2_weights[58][76] = 16'sd23;
        fc2_weights[58][77] = 16'sd-9;
        fc2_weights[58][78] = 16'sd-1;
        fc2_weights[58][79] = 16'sd-17;
        fc2_weights[58][80] = 16'sd-59;
        fc2_weights[58][81] = 16'sd15;
        fc2_weights[58][82] = 16'sd-37;
        fc2_weights[58][83] = 16'sd5;
        fc2_weights[58][84] = 16'sd-3;
        fc2_weights[58][85] = 16'sd-25;
        fc2_weights[58][86] = 16'sd-24;
        fc2_weights[58][87] = 16'sd-46;
        fc2_weights[58][88] = 16'sd1;
        fc2_weights[58][89] = 16'sd-35;
        fc2_weights[58][90] = 16'sd-18;
        fc2_weights[58][91] = 16'sd2;
        fc2_weights[58][92] = 16'sd-9;
        fc2_weights[58][93] = 16'sd-25;
        fc2_weights[58][94] = 16'sd18;
        fc2_weights[58][95] = 16'sd-8;
        fc2_weights[58][96] = 16'sd34;
        fc2_weights[58][97] = 16'sd-22;
        fc2_weights[58][98] = 16'sd-16;
        fc2_weights[58][99] = 16'sd-89;
        fc2_weights[58][100] = 16'sd51;
        fc2_weights[58][101] = 16'sd-55;
        fc2_weights[58][102] = 16'sd5;
        fc2_weights[58][103] = 16'sd74;
        fc2_weights[58][104] = 16'sd103;
        fc2_weights[58][105] = 16'sd-10;
        fc2_weights[58][106] = 16'sd-25;
        fc2_weights[58][107] = 16'sd-33;
        fc2_weights[58][108] = 16'sd-53;
        fc2_weights[58][109] = 16'sd14;
        fc2_weights[58][110] = 16'sd5;
        fc2_weights[58][111] = 16'sd-26;
        fc2_weights[58][112] = 16'sd-39;
        fc2_weights[58][113] = 16'sd-53;
        fc2_weights[58][114] = 16'sd9;
        fc2_weights[58][115] = 16'sd-46;
        fc2_weights[58][116] = 16'sd15;
        fc2_weights[58][117] = 16'sd58;
        fc2_weights[58][118] = 16'sd-67;
        fc2_weights[58][119] = 16'sd-20;
        fc2_weights[58][120] = 16'sd-52;
        fc2_weights[58][121] = 16'sd-60;
        fc2_weights[58][122] = 16'sd-2;
        fc2_weights[58][123] = 16'sd20;
        fc2_weights[58][124] = 16'sd-41;
        fc2_weights[58][125] = 16'sd4;
        fc2_weights[58][126] = 16'sd-14;
        fc2_weights[58][127] = 16'sd48;
        fc2_weights[59][0] = 16'sd-41;
        fc2_weights[59][1] = 16'sd-9;
        fc2_weights[59][2] = 16'sd45;
        fc2_weights[59][3] = 16'sd-4;
        fc2_weights[59][4] = 16'sd-38;
        fc2_weights[59][5] = 16'sd-44;
        fc2_weights[59][6] = 16'sd-30;
        fc2_weights[59][7] = 16'sd-39;
        fc2_weights[59][8] = 16'sd-51;
        fc2_weights[59][9] = 16'sd25;
        fc2_weights[59][10] = 16'sd-49;
        fc2_weights[59][11] = 16'sd-53;
        fc2_weights[59][12] = 16'sd-7;
        fc2_weights[59][13] = 16'sd24;
        fc2_weights[59][14] = 16'sd2;
        fc2_weights[59][15] = 16'sd54;
        fc2_weights[59][16] = 16'sd-28;
        fc2_weights[59][17] = 16'sd12;
        fc2_weights[59][18] = 16'sd25;
        fc2_weights[59][19] = 16'sd14;
        fc2_weights[59][20] = 16'sd-6;
        fc2_weights[59][21] = 16'sd6;
        fc2_weights[59][22] = 16'sd-23;
        fc2_weights[59][23] = 16'sd28;
        fc2_weights[59][24] = 16'sd26;
        fc2_weights[59][25] = 16'sd-20;
        fc2_weights[59][26] = 16'sd-63;
        fc2_weights[59][27] = 16'sd-22;
        fc2_weights[59][28] = 16'sd-35;
        fc2_weights[59][29] = 16'sd-17;
        fc2_weights[59][30] = 16'sd-18;
        fc2_weights[59][31] = 16'sd-58;
        fc2_weights[59][32] = 16'sd29;
        fc2_weights[59][33] = 16'sd-24;
        fc2_weights[59][34] = 16'sd49;
        fc2_weights[59][35] = 16'sd-21;
        fc2_weights[59][36] = 16'sd-24;
        fc2_weights[59][37] = 16'sd0;
        fc2_weights[59][38] = 16'sd-76;
        fc2_weights[59][39] = 16'sd-39;
        fc2_weights[59][40] = 16'sd23;
        fc2_weights[59][41] = 16'sd23;
        fc2_weights[59][42] = 16'sd-44;
        fc2_weights[59][43] = 16'sd7;
        fc2_weights[59][44] = 16'sd51;
        fc2_weights[59][45] = 16'sd43;
        fc2_weights[59][46] = 16'sd14;
        fc2_weights[59][47] = 16'sd-13;
        fc2_weights[59][48] = 16'sd-8;
        fc2_weights[59][49] = 16'sd16;
        fc2_weights[59][50] = 16'sd-8;
        fc2_weights[59][51] = 16'sd-7;
        fc2_weights[59][52] = 16'sd102;
        fc2_weights[59][53] = 16'sd-20;
        fc2_weights[59][54] = 16'sd19;
        fc2_weights[59][55] = 16'sd-12;
        fc2_weights[59][56] = 16'sd-42;
        fc2_weights[59][57] = 16'sd8;
        fc2_weights[59][58] = 16'sd-33;
        fc2_weights[59][59] = 16'sd51;
        fc2_weights[59][60] = 16'sd32;
        fc2_weights[59][61] = 16'sd-76;
        fc2_weights[59][62] = 16'sd-26;
        fc2_weights[59][63] = 16'sd71;
        fc2_weights[59][64] = 16'sd-32;
        fc2_weights[59][65] = 16'sd66;
        fc2_weights[59][66] = 16'sd37;
        fc2_weights[59][67] = 16'sd-57;
        fc2_weights[59][68] = 16'sd63;
        fc2_weights[59][69] = 16'sd59;
        fc2_weights[59][70] = 16'sd-12;
        fc2_weights[59][71] = 16'sd-37;
        fc2_weights[59][72] = 16'sd-4;
        fc2_weights[59][73] = 16'sd-22;
        fc2_weights[59][74] = 16'sd2;
        fc2_weights[59][75] = 16'sd-8;
        fc2_weights[59][76] = 16'sd23;
        fc2_weights[59][77] = 16'sd-48;
        fc2_weights[59][78] = 16'sd-20;
        fc2_weights[59][79] = 16'sd-2;
        fc2_weights[59][80] = 16'sd-74;
        fc2_weights[59][81] = 16'sd-63;
        fc2_weights[59][82] = 16'sd-90;
        fc2_weights[59][83] = 16'sd-12;
        fc2_weights[59][84] = 16'sd46;
        fc2_weights[59][85] = 16'sd-42;
        fc2_weights[59][86] = 16'sd27;
        fc2_weights[59][87] = 16'sd-64;
        fc2_weights[59][88] = 16'sd66;
        fc2_weights[59][89] = 16'sd-18;
        fc2_weights[59][90] = 16'sd79;
        fc2_weights[59][91] = 16'sd-12;
        fc2_weights[59][92] = 16'sd64;
        fc2_weights[59][93] = 16'sd-47;
        fc2_weights[59][94] = 16'sd-8;
        fc2_weights[59][95] = 16'sd-29;
        fc2_weights[59][96] = 16'sd-12;
        fc2_weights[59][97] = 16'sd-29;
        fc2_weights[59][98] = 16'sd-33;
        fc2_weights[59][99] = 16'sd-41;
        fc2_weights[59][100] = 16'sd32;
        fc2_weights[59][101] = 16'sd25;
        fc2_weights[59][102] = 16'sd-22;
        fc2_weights[59][103] = 16'sd-34;
        fc2_weights[59][104] = 16'sd64;
        fc2_weights[59][105] = 16'sd-61;
        fc2_weights[59][106] = 16'sd-71;
        fc2_weights[59][107] = 16'sd19;
        fc2_weights[59][108] = 16'sd-25;
        fc2_weights[59][109] = 16'sd-21;
        fc2_weights[59][110] = 16'sd10;
        fc2_weights[59][111] = 16'sd14;
        fc2_weights[59][112] = 16'sd-42;
        fc2_weights[59][113] = 16'sd-58;
        fc2_weights[59][114] = 16'sd-11;
        fc2_weights[59][115] = 16'sd-24;
        fc2_weights[59][116] = 16'sd40;
        fc2_weights[59][117] = 16'sd44;
        fc2_weights[59][118] = 16'sd-49;
        fc2_weights[59][119] = 16'sd-65;
        fc2_weights[59][120] = 16'sd-56;
        fc2_weights[59][121] = 16'sd-10;
        fc2_weights[59][122] = 16'sd46;
        fc2_weights[59][123] = 16'sd0;
        fc2_weights[59][124] = 16'sd-27;
        fc2_weights[59][125] = 16'sd45;
        fc2_weights[59][126] = 16'sd10;
        fc2_weights[59][127] = 16'sd74;
        fc2_weights[60][0] = 16'sd82;
        fc2_weights[60][1] = 16'sd-1;
        fc2_weights[60][2] = 16'sd30;
        fc2_weights[60][3] = 16'sd48;
        fc2_weights[60][4] = 16'sd36;
        fc2_weights[60][5] = 16'sd53;
        fc2_weights[60][6] = 16'sd56;
        fc2_weights[60][7] = 16'sd-56;
        fc2_weights[60][8] = 16'sd23;
        fc2_weights[60][9] = 16'sd21;
        fc2_weights[60][10] = 16'sd-9;
        fc2_weights[60][11] = 16'sd17;
        fc2_weights[60][12] = 16'sd-56;
        fc2_weights[60][13] = 16'sd44;
        fc2_weights[60][14] = 16'sd8;
        fc2_weights[60][15] = 16'sd4;
        fc2_weights[60][16] = 16'sd37;
        fc2_weights[60][17] = 16'sd-54;
        fc2_weights[60][18] = 16'sd15;
        fc2_weights[60][19] = 16'sd36;
        fc2_weights[60][20] = 16'sd-33;
        fc2_weights[60][21] = 16'sd-28;
        fc2_weights[60][22] = 16'sd-9;
        fc2_weights[60][23] = 16'sd38;
        fc2_weights[60][24] = 16'sd10;
        fc2_weights[60][25] = 16'sd-23;
        fc2_weights[60][26] = 16'sd-19;
        fc2_weights[60][27] = 16'sd-15;
        fc2_weights[60][28] = 16'sd25;
        fc2_weights[60][29] = 16'sd30;
        fc2_weights[60][30] = 16'sd2;
        fc2_weights[60][31] = 16'sd49;
        fc2_weights[60][32] = 16'sd-40;
        fc2_weights[60][33] = 16'sd13;
        fc2_weights[60][34] = 16'sd9;
        fc2_weights[60][35] = 16'sd26;
        fc2_weights[60][36] = 16'sd-16;
        fc2_weights[60][37] = 16'sd-74;
        fc2_weights[60][38] = 16'sd41;
        fc2_weights[60][39] = 16'sd12;
        fc2_weights[60][40] = 16'sd16;
        fc2_weights[60][41] = 16'sd46;
        fc2_weights[60][42] = 16'sd-25;
        fc2_weights[60][43] = 16'sd3;
        fc2_weights[60][44] = 16'sd-15;
        fc2_weights[60][45] = 16'sd-19;
        fc2_weights[60][46] = 16'sd30;
        fc2_weights[60][47] = 16'sd1;
        fc2_weights[60][48] = 16'sd16;
        fc2_weights[60][49] = 16'sd21;
        fc2_weights[60][50] = 16'sd-23;
        fc2_weights[60][51] = 16'sd9;
        fc2_weights[60][52] = 16'sd18;
        fc2_weights[60][53] = 16'sd41;
        fc2_weights[60][54] = 16'sd-15;
        fc2_weights[60][55] = 16'sd64;
        fc2_weights[60][56] = 16'sd-9;
        fc2_weights[60][57] = 16'sd17;
        fc2_weights[60][58] = 16'sd7;
        fc2_weights[60][59] = 16'sd-47;
        fc2_weights[60][60] = 16'sd22;
        fc2_weights[60][61] = 16'sd10;
        fc2_weights[60][62] = 16'sd74;
        fc2_weights[60][63] = 16'sd-3;
        fc2_weights[60][64] = 16'sd9;
        fc2_weights[60][65] = 16'sd23;
        fc2_weights[60][66] = 16'sd58;
        fc2_weights[60][67] = 16'sd-40;
        fc2_weights[60][68] = 16'sd0;
        fc2_weights[60][69] = 16'sd-61;
        fc2_weights[60][70] = 16'sd-13;
        fc2_weights[60][71] = 16'sd22;
        fc2_weights[60][72] = 16'sd7;
        fc2_weights[60][73] = 16'sd20;
        fc2_weights[60][74] = 16'sd-21;
        fc2_weights[60][75] = 16'sd-1;
        fc2_weights[60][76] = 16'sd4;
        fc2_weights[60][77] = 16'sd28;
        fc2_weights[60][78] = 16'sd-36;
        fc2_weights[60][79] = 16'sd6;
        fc2_weights[60][80] = 16'sd42;
        fc2_weights[60][81] = 16'sd12;
        fc2_weights[60][82] = 16'sd-30;
        fc2_weights[60][83] = 16'sd26;
        fc2_weights[60][84] = 16'sd19;
        fc2_weights[60][85] = 16'sd44;
        fc2_weights[60][86] = 16'sd12;
        fc2_weights[60][87] = 16'sd-4;
        fc2_weights[60][88] = 16'sd-3;
        fc2_weights[60][89] = 16'sd53;
        fc2_weights[60][90] = 16'sd5;
        fc2_weights[60][91] = 16'sd4;
        fc2_weights[60][92] = 16'sd67;
        fc2_weights[60][93] = 16'sd17;
        fc2_weights[60][94] = 16'sd-110;
        fc2_weights[60][95] = 16'sd-48;
        fc2_weights[60][96] = 16'sd-55;
        fc2_weights[60][97] = 16'sd14;
        fc2_weights[60][98] = 16'sd18;
        fc2_weights[60][99] = 16'sd-10;
        fc2_weights[60][100] = 16'sd10;
        fc2_weights[60][101] = 16'sd26;
        fc2_weights[60][102] = 16'sd-4;
        fc2_weights[60][103] = 16'sd-15;
        fc2_weights[60][104] = 16'sd64;
        fc2_weights[60][105] = 16'sd8;
        fc2_weights[60][106] = 16'sd-25;
        fc2_weights[60][107] = 16'sd64;
        fc2_weights[60][108] = 16'sd-59;
        fc2_weights[60][109] = 16'sd27;
        fc2_weights[60][110] = 16'sd3;
        fc2_weights[60][111] = 16'sd-31;
        fc2_weights[60][112] = 16'sd4;
        fc2_weights[60][113] = 16'sd18;
        fc2_weights[60][114] = 16'sd63;
        fc2_weights[60][115] = 16'sd44;
        fc2_weights[60][116] = 16'sd-28;
        fc2_weights[60][117] = 16'sd-33;
        fc2_weights[60][118] = 16'sd41;
        fc2_weights[60][119] = 16'sd78;
        fc2_weights[60][120] = 16'sd-21;
        fc2_weights[60][121] = 16'sd-11;
        fc2_weights[60][122] = 16'sd-10;
        fc2_weights[60][123] = 16'sd22;
        fc2_weights[60][124] = 16'sd-15;
        fc2_weights[60][125] = 16'sd-37;
        fc2_weights[60][126] = 16'sd4;
        fc2_weights[60][127] = 16'sd-18;
        fc2_weights[61][0] = 16'sd-1;
        fc2_weights[61][1] = 16'sd-36;
        fc2_weights[61][2] = 16'sd50;
        fc2_weights[61][3] = 16'sd9;
        fc2_weights[61][4] = 16'sd-29;
        fc2_weights[61][5] = 16'sd3;
        fc2_weights[61][6] = 16'sd-6;
        fc2_weights[61][7] = 16'sd-9;
        fc2_weights[61][8] = 16'sd-17;
        fc2_weights[61][9] = 16'sd30;
        fc2_weights[61][10] = 16'sd-21;
        fc2_weights[61][11] = 16'sd-18;
        fc2_weights[61][12] = 16'sd8;
        fc2_weights[61][13] = 16'sd35;
        fc2_weights[61][14] = 16'sd61;
        fc2_weights[61][15] = 16'sd22;
        fc2_weights[61][16] = 16'sd2;
        fc2_weights[61][17] = 16'sd70;
        fc2_weights[61][18] = 16'sd129;
        fc2_weights[61][19] = 16'sd-19;
        fc2_weights[61][20] = 16'sd48;
        fc2_weights[61][21] = 16'sd-25;
        fc2_weights[61][22] = 16'sd7;
        fc2_weights[61][23] = 16'sd-7;
        fc2_weights[61][24] = 16'sd-4;
        fc2_weights[61][25] = 16'sd12;
        fc2_weights[61][26] = 16'sd-54;
        fc2_weights[61][27] = 16'sd22;
        fc2_weights[61][28] = 16'sd-58;
        fc2_weights[61][29] = 16'sd-29;
        fc2_weights[61][30] = 16'sd37;
        fc2_weights[61][31] = 16'sd-14;
        fc2_weights[61][32] = 16'sd-29;
        fc2_weights[61][33] = 16'sd-4;
        fc2_weights[61][34] = 16'sd4;
        fc2_weights[61][35] = 16'sd-37;
        fc2_weights[61][36] = 16'sd-14;
        fc2_weights[61][37] = 16'sd5;
        fc2_weights[61][38] = 16'sd-58;
        fc2_weights[61][39] = 16'sd-59;
        fc2_weights[61][40] = 16'sd-5;
        fc2_weights[61][41] = 16'sd42;
        fc2_weights[61][42] = 16'sd22;
        fc2_weights[61][43] = 16'sd25;
        fc2_weights[61][44] = 16'sd-4;
        fc2_weights[61][45] = 16'sd-32;
        fc2_weights[61][46] = 16'sd39;
        fc2_weights[61][47] = 16'sd-36;
        fc2_weights[61][48] = 16'sd47;
        fc2_weights[61][49] = 16'sd4;
        fc2_weights[61][50] = 16'sd45;
        fc2_weights[61][51] = 16'sd3;
        fc2_weights[61][52] = 16'sd139;
        fc2_weights[61][53] = 16'sd-6;
        fc2_weights[61][54] = 16'sd18;
        fc2_weights[61][55] = 16'sd-9;
        fc2_weights[61][56] = 16'sd24;
        fc2_weights[61][57] = 16'sd-26;
        fc2_weights[61][58] = 16'sd55;
        fc2_weights[61][59] = 16'sd29;
        fc2_weights[61][60] = 16'sd-4;
        fc2_weights[61][61] = 16'sd-65;
        fc2_weights[61][62] = 16'sd38;
        fc2_weights[61][63] = 16'sd17;
        fc2_weights[61][64] = 16'sd-15;
        fc2_weights[61][65] = 16'sd63;
        fc2_weights[61][66] = 16'sd-8;
        fc2_weights[61][67] = 16'sd28;
        fc2_weights[61][68] = 16'sd-32;
        fc2_weights[61][69] = 16'sd6;
        fc2_weights[61][70] = 16'sd-5;
        fc2_weights[61][71] = 16'sd-59;
        fc2_weights[61][72] = 16'sd68;
        fc2_weights[61][73] = 16'sd-4;
        fc2_weights[61][74] = 16'sd-4;
        fc2_weights[61][75] = 16'sd-30;
        fc2_weights[61][76] = 16'sd-68;
        fc2_weights[61][77] = 16'sd-12;
        fc2_weights[61][78] = 16'sd-18;
        fc2_weights[61][79] = 16'sd-8;
        fc2_weights[61][80] = 16'sd-37;
        fc2_weights[61][81] = 16'sd44;
        fc2_weights[61][82] = 16'sd-1;
        fc2_weights[61][83] = 16'sd-10;
        fc2_weights[61][84] = 16'sd-5;
        fc2_weights[61][85] = 16'sd-22;
        fc2_weights[61][86] = 16'sd-45;
        fc2_weights[61][87] = 16'sd-52;
        fc2_weights[61][88] = 16'sd38;
        fc2_weights[61][89] = 16'sd4;
        fc2_weights[61][90] = 16'sd12;
        fc2_weights[61][91] = 16'sd-13;
        fc2_weights[61][92] = 16'sd16;
        fc2_weights[61][93] = 16'sd-37;
        fc2_weights[61][94] = 16'sd55;
        fc2_weights[61][95] = 16'sd-19;
        fc2_weights[61][96] = 16'sd-21;
        fc2_weights[61][97] = 16'sd2;
        fc2_weights[61][98] = 16'sd-36;
        fc2_weights[61][99] = 16'sd-9;
        fc2_weights[61][100] = 16'sd-14;
        fc2_weights[61][101] = 16'sd5;
        fc2_weights[61][102] = 16'sd18;
        fc2_weights[61][103] = 16'sd46;
        fc2_weights[61][104] = 16'sd-1;
        fc2_weights[61][105] = 16'sd-2;
        fc2_weights[61][106] = 16'sd-3;
        fc2_weights[61][107] = 16'sd28;
        fc2_weights[61][108] = 16'sd35;
        fc2_weights[61][109] = 16'sd-21;
        fc2_weights[61][110] = 16'sd43;
        fc2_weights[61][111] = 16'sd-2;
        fc2_weights[61][112] = 16'sd-27;
        fc2_weights[61][113] = 16'sd-59;
        fc2_weights[61][114] = 16'sd-3;
        fc2_weights[61][115] = 16'sd-18;
        fc2_weights[61][116] = 16'sd17;
        fc2_weights[61][117] = 16'sd7;
        fc2_weights[61][118] = 16'sd10;
        fc2_weights[61][119] = 16'sd-11;
        fc2_weights[61][120] = 16'sd11;
        fc2_weights[61][121] = 16'sd16;
        fc2_weights[61][122] = 16'sd54;
        fc2_weights[61][123] = 16'sd21;
        fc2_weights[61][124] = 16'sd-22;
        fc2_weights[61][125] = 16'sd22;
        fc2_weights[61][126] = 16'sd22;
        fc2_weights[61][127] = 16'sd-27;
        fc2_weights[62][0] = 16'sd22;
        fc2_weights[62][1] = 16'sd43;
        fc2_weights[62][2] = 16'sd48;
        fc2_weights[62][3] = 16'sd4;
        fc2_weights[62][4] = 16'sd9;
        fc2_weights[62][5] = 16'sd-18;
        fc2_weights[62][6] = 16'sd-5;
        fc2_weights[62][7] = 16'sd-20;
        fc2_weights[62][8] = 16'sd55;
        fc2_weights[62][9] = 16'sd8;
        fc2_weights[62][10] = 16'sd-39;
        fc2_weights[62][11] = 16'sd38;
        fc2_weights[62][12] = 16'sd0;
        fc2_weights[62][13] = 16'sd-4;
        fc2_weights[62][14] = 16'sd-19;
        fc2_weights[62][15] = 16'sd-8;
        fc2_weights[62][16] = 16'sd-3;
        fc2_weights[62][17] = 16'sd-29;
        fc2_weights[62][18] = 16'sd-49;
        fc2_weights[62][19] = 16'sd-34;
        fc2_weights[62][20] = 16'sd-37;
        fc2_weights[62][21] = 16'sd-33;
        fc2_weights[62][22] = 16'sd-64;
        fc2_weights[62][23] = 16'sd22;
        fc2_weights[62][24] = 16'sd-14;
        fc2_weights[62][25] = 16'sd-36;
        fc2_weights[62][26] = 16'sd-6;
        fc2_weights[62][27] = 16'sd-41;
        fc2_weights[62][28] = 16'sd79;
        fc2_weights[62][29] = 16'sd-24;
        fc2_weights[62][30] = 16'sd26;
        fc2_weights[62][31] = 16'sd62;
        fc2_weights[62][32] = 16'sd18;
        fc2_weights[62][33] = 16'sd-21;
        fc2_weights[62][34] = 16'sd-28;
        fc2_weights[62][35] = 16'sd-34;
        fc2_weights[62][36] = 16'sd-32;
        fc2_weights[62][37] = 16'sd1;
        fc2_weights[62][38] = 16'sd31;
        fc2_weights[62][39] = 16'sd54;
        fc2_weights[62][40] = 16'sd-12;
        fc2_weights[62][41] = 16'sd-18;
        fc2_weights[62][42] = 16'sd16;
        fc2_weights[62][43] = 16'sd4;
        fc2_weights[62][44] = 16'sd-57;
        fc2_weights[62][45] = 16'sd-102;
        fc2_weights[62][46] = 16'sd6;
        fc2_weights[62][47] = 16'sd86;
        fc2_weights[62][48] = 16'sd-5;
        fc2_weights[62][49] = 16'sd2;
        fc2_weights[62][50] = 16'sd-23;
        fc2_weights[62][51] = 16'sd-26;
        fc2_weights[62][52] = 16'sd-38;
        fc2_weights[62][53] = 16'sd-19;
        fc2_weights[62][54] = 16'sd-7;
        fc2_weights[62][55] = 16'sd61;
        fc2_weights[62][56] = 16'sd41;
        fc2_weights[62][57] = 16'sd-2;
        fc2_weights[62][58] = 16'sd-54;
        fc2_weights[62][59] = 16'sd-7;
        fc2_weights[62][60] = 16'sd-74;
        fc2_weights[62][61] = 16'sd-13;
        fc2_weights[62][62] = 16'sd-35;
        fc2_weights[62][63] = 16'sd-30;
        fc2_weights[62][64] = 16'sd40;
        fc2_weights[62][65] = 16'sd-39;
        fc2_weights[62][66] = 16'sd-68;
        fc2_weights[62][67] = 16'sd-22;
        fc2_weights[62][68] = 16'sd-51;
        fc2_weights[62][69] = 16'sd6;
        fc2_weights[62][70] = 16'sd40;
        fc2_weights[62][71] = 16'sd-45;
        fc2_weights[62][72] = 16'sd68;
        fc2_weights[62][73] = 16'sd20;
        fc2_weights[62][74] = 16'sd-32;
        fc2_weights[62][75] = 16'sd-17;
        fc2_weights[62][76] = 16'sd-17;
        fc2_weights[62][77] = 16'sd-35;
        fc2_weights[62][78] = 16'sd-42;
        fc2_weights[62][79] = 16'sd22;
        fc2_weights[62][80] = 16'sd81;
        fc2_weights[62][81] = 16'sd-62;
        fc2_weights[62][82] = 16'sd-39;
        fc2_weights[62][83] = 16'sd43;
        fc2_weights[62][84] = 16'sd40;
        fc2_weights[62][85] = 16'sd17;
        fc2_weights[62][86] = 16'sd31;
        fc2_weights[62][87] = 16'sd-48;
        fc2_weights[62][88] = 16'sd-33;
        fc2_weights[62][89] = 16'sd27;
        fc2_weights[62][90] = 16'sd-71;
        fc2_weights[62][91] = 16'sd-17;
        fc2_weights[62][92] = 16'sd-40;
        fc2_weights[62][93] = 16'sd32;
        fc2_weights[62][94] = 16'sd-8;
        fc2_weights[62][95] = 16'sd-19;
        fc2_weights[62][96] = 16'sd3;
        fc2_weights[62][97] = 16'sd-5;
        fc2_weights[62][98] = 16'sd56;
        fc2_weights[62][99] = 16'sd-22;
        fc2_weights[62][100] = 16'sd-60;
        fc2_weights[62][101] = 16'sd10;
        fc2_weights[62][102] = 16'sd-9;
        fc2_weights[62][103] = 16'sd-29;
        fc2_weights[62][104] = 16'sd26;
        fc2_weights[62][105] = 16'sd0;
        fc2_weights[62][106] = 16'sd-28;
        fc2_weights[62][107] = 16'sd24;
        fc2_weights[62][108] = 16'sd-30;
        fc2_weights[62][109] = 16'sd1;
        fc2_weights[62][110] = 16'sd-59;
        fc2_weights[62][111] = 16'sd-60;
        fc2_weights[62][112] = 16'sd75;
        fc2_weights[62][113] = 16'sd8;
        fc2_weights[62][114] = 16'sd-66;
        fc2_weights[62][115] = 16'sd-9;
        fc2_weights[62][116] = 16'sd-42;
        fc2_weights[62][117] = 16'sd-15;
        fc2_weights[62][118] = 16'sd9;
        fc2_weights[62][119] = 16'sd21;
        fc2_weights[62][120] = 16'sd-17;
        fc2_weights[62][121] = 16'sd-33;
        fc2_weights[62][122] = 16'sd-73;
        fc2_weights[62][123] = 16'sd13;
        fc2_weights[62][124] = 16'sd0;
        fc2_weights[62][125] = 16'sd6;
        fc2_weights[62][126] = 16'sd-38;
        fc2_weights[62][127] = 16'sd-80;
        fc2_weights[63][0] = 16'sd30;
        fc2_weights[63][1] = 16'sd19;
        fc2_weights[63][2] = 16'sd19;
        fc2_weights[63][3] = 16'sd37;
        fc2_weights[63][4] = 16'sd-5;
        fc2_weights[63][5] = 16'sd-37;
        fc2_weights[63][6] = 16'sd55;
        fc2_weights[63][7] = 16'sd-11;
        fc2_weights[63][8] = 16'sd120;
        fc2_weights[63][9] = 16'sd-20;
        fc2_weights[63][10] = 16'sd-28;
        fc2_weights[63][11] = 16'sd-15;
        fc2_weights[63][12] = 16'sd61;
        fc2_weights[63][13] = 16'sd-14;
        fc2_weights[63][14] = 16'sd-70;
        fc2_weights[63][15] = 16'sd0;
        fc2_weights[63][16] = 16'sd-30;
        fc2_weights[63][17] = 16'sd54;
        fc2_weights[63][18] = 16'sd-19;
        fc2_weights[63][19] = 16'sd-56;
        fc2_weights[63][20] = 16'sd43;
        fc2_weights[63][21] = 16'sd-16;
        fc2_weights[63][22] = 16'sd-35;
        fc2_weights[63][23] = 16'sd-7;
        fc2_weights[63][24] = 16'sd-22;
        fc2_weights[63][25] = 16'sd-9;
        fc2_weights[63][26] = 16'sd-19;
        fc2_weights[63][27] = 16'sd-23;
        fc2_weights[63][28] = 16'sd40;
        fc2_weights[63][29] = 16'sd27;
        fc2_weights[63][30] = 16'sd6;
        fc2_weights[63][31] = 16'sd15;
        fc2_weights[63][32] = 16'sd55;
        fc2_weights[63][33] = 16'sd40;
        fc2_weights[63][34] = 16'sd-6;
        fc2_weights[63][35] = 16'sd7;
        fc2_weights[63][36] = 16'sd-23;
        fc2_weights[63][37] = 16'sd-36;
        fc2_weights[63][38] = 16'sd10;
        fc2_weights[63][39] = 16'sd35;
        fc2_weights[63][40] = 16'sd-47;
        fc2_weights[63][41] = 16'sd-30;
        fc2_weights[63][42] = 16'sd73;
        fc2_weights[63][43] = 16'sd33;
        fc2_weights[63][44] = 16'sd-30;
        fc2_weights[63][45] = 16'sd-39;
        fc2_weights[63][46] = 16'sd-36;
        fc2_weights[63][47] = 16'sd37;
        fc2_weights[63][48] = 16'sd23;
        fc2_weights[63][49] = 16'sd-72;
        fc2_weights[63][50] = 16'sd5;
        fc2_weights[63][51] = 16'sd-80;
        fc2_weights[63][52] = 16'sd-11;
        fc2_weights[63][53] = 16'sd-34;
        fc2_weights[63][54] = 16'sd-23;
        fc2_weights[63][55] = 16'sd32;
        fc2_weights[63][56] = 16'sd49;
        fc2_weights[63][57] = 16'sd-78;
        fc2_weights[63][58] = 16'sd4;
        fc2_weights[63][59] = 16'sd-36;
        fc2_weights[63][60] = 16'sd-32;
        fc2_weights[63][61] = 16'sd25;
        fc2_weights[63][62] = 16'sd-91;
        fc2_weights[63][63] = 16'sd-56;
        fc2_weights[63][64] = 16'sd-19;
        fc2_weights[63][65] = 16'sd23;
        fc2_weights[63][66] = 16'sd-101;
        fc2_weights[63][67] = 16'sd2;
        fc2_weights[63][68] = 16'sd-8;
        fc2_weights[63][69] = 16'sd-21;
        fc2_weights[63][70] = 16'sd-13;
        fc2_weights[63][71] = 16'sd-34;
        fc2_weights[63][72] = 16'sd22;
        fc2_weights[63][73] = 16'sd-9;
        fc2_weights[63][74] = 16'sd-24;
        fc2_weights[63][75] = 16'sd-7;
        fc2_weights[63][76] = 16'sd-14;
        fc2_weights[63][77] = 16'sd-41;
        fc2_weights[63][78] = 16'sd10;
        fc2_weights[63][79] = 16'sd-9;
        fc2_weights[63][80] = 16'sd-32;
        fc2_weights[63][81] = 16'sd-74;
        fc2_weights[63][82] = 16'sd-4;
        fc2_weights[63][83] = 16'sd-22;
        fc2_weights[63][84] = 16'sd-2;
        fc2_weights[63][85] = 16'sd18;
        fc2_weights[63][86] = 16'sd-15;
        fc2_weights[63][87] = 16'sd-42;
        fc2_weights[63][88] = 16'sd-4;
        fc2_weights[63][89] = 16'sd-13;
        fc2_weights[63][90] = 16'sd-30;
        fc2_weights[63][91] = 16'sd-31;
        fc2_weights[63][92] = 16'sd-55;
        fc2_weights[63][93] = 16'sd119;
        fc2_weights[63][94] = 16'sd-38;
        fc2_weights[63][95] = 16'sd-57;
        fc2_weights[63][96] = 16'sd29;
        fc2_weights[63][97] = 16'sd13;
        fc2_weights[63][98] = 16'sd-5;
        fc2_weights[63][99] = 16'sd-2;
        fc2_weights[63][100] = 16'sd-73;
        fc2_weights[63][101] = 16'sd-26;
        fc2_weights[63][102] = 16'sd-60;
        fc2_weights[63][103] = 16'sd-91;
        fc2_weights[63][104] = 16'sd-8;
        fc2_weights[63][105] = 16'sd13;
        fc2_weights[63][106] = 16'sd-57;
        fc2_weights[63][107] = 16'sd10;
        fc2_weights[63][108] = 16'sd-46;
        fc2_weights[63][109] = 16'sd-6;
        fc2_weights[63][110] = 16'sd-72;
        fc2_weights[63][111] = 16'sd-55;
        fc2_weights[63][112] = 16'sd54;
        fc2_weights[63][113] = 16'sd88;
        fc2_weights[63][114] = 16'sd-62;
        fc2_weights[63][115] = 16'sd-14;
        fc2_weights[63][116] = 16'sd-10;
        fc2_weights[63][117] = 16'sd62;
        fc2_weights[63][118] = 16'sd18;
        fc2_weights[63][119] = 16'sd54;
        fc2_weights[63][120] = 16'sd4;
        fc2_weights[63][121] = 16'sd-1;
        fc2_weights[63][122] = 16'sd-54;
        fc2_weights[63][123] = 16'sd-25;
        fc2_weights[63][124] = 16'sd-28;
        fc2_weights[63][125] = 16'sd-35;
        fc2_weights[63][126] = 16'sd-62;
        fc2_weights[63][127] = 16'sd-30;
        // fc2 biases
        fc2_biases[0] = 16'sd0;
        fc2_biases[1] = 16'sd0;
        fc2_biases[2] = 16'sd0;
        fc2_biases[3] = 16'sd0;
        fc2_biases[4] = 16'sd0;
        fc2_biases[5] = 16'sd0;
        fc2_biases[6] = 16'sd0;
        fc2_biases[7] = 16'sd0;
        fc2_biases[8] = 16'sd0;
        fc2_biases[9] = 16'sd0;
        fc2_biases[10] = 16'sd0;
        fc2_biases[11] = 16'sd0;
        fc2_biases[12] = 16'sd0;
        fc2_biases[13] = 16'sd0;
        fc2_biases[14] = 16'sd0;
        fc2_biases[15] = 16'sd0;
        fc2_biases[16] = 16'sd0;
        fc2_biases[17] = 16'sd0;
        fc2_biases[18] = 16'sd0;
        fc2_biases[19] = 16'sd0;
        fc2_biases[20] = 16'sd0;
        fc2_biases[21] = 16'sd0;
        fc2_biases[22] = 16'sd0;
        fc2_biases[23] = 16'sd0;
        fc2_biases[24] = 16'sd0;
        fc2_biases[25] = 16'sd0;
        fc2_biases[26] = 16'sd0;
        fc2_biases[27] = 16'sd0;
        fc2_biases[28] = 16'sd0;
        fc2_biases[29] = 16'sd0;
        fc2_biases[30] = 16'sd0;
        fc2_biases[31] = 16'sd0;
        fc2_biases[32] = 16'sd0;
        fc2_biases[33] = 16'sd0;
        fc2_biases[34] = 16'sd0;
        fc2_biases[35] = 16'sd0;
        fc2_biases[36] = 16'sd0;
        fc2_biases[37] = 16'sd0;
        fc2_biases[38] = 16'sd0;
        fc2_biases[39] = 16'sd0;
        fc2_biases[40] = 16'sd0;
        fc2_biases[41] = 16'sd0;
        fc2_biases[42] = 16'sd0;
        fc2_biases[43] = 16'sd0;
        fc2_biases[44] = 16'sd0;
        fc2_biases[45] = 16'sd0;
        fc2_biases[46] = 16'sd0;
        fc2_biases[47] = 16'sd0;
        fc2_biases[48] = 16'sd0;
        fc2_biases[49] = 16'sd0;
        fc2_biases[50] = 16'sd0;
        fc2_biases[51] = 16'sd0;
        fc2_biases[52] = 16'sd0;
        fc2_biases[53] = 16'sd0;
        fc2_biases[54] = 16'sd0;
        fc2_biases[55] = 16'sd0;
        fc2_biases[56] = 16'sd0;
        fc2_biases[57] = 16'sd0;
        fc2_biases[58] = 16'sd0;
        fc2_biases[59] = 16'sd0;
        fc2_biases[60] = 16'sd0;
        fc2_biases[61] = 16'sd0;
        fc2_biases[62] = 16'sd0;
        fc2_biases[63] = 16'sd0;
        
        // fc3 weights
        fc3_weights[0][0] = 16'sd1;
        fc3_weights[0][1] = 16'sd-7;
        fc3_weights[0][2] = 16'sd0;
        fc3_weights[0][3] = 16'sd-4;
        fc3_weights[0][4] = 16'sd14;
        fc3_weights[0][5] = 16'sd-1;
        fc3_weights[0][6] = 16'sd34;
        fc3_weights[0][7] = 16'sd-15;
        fc3_weights[0][8] = 16'sd-2;
        fc3_weights[0][9] = 16'sd12;
        fc3_weights[0][10] = 16'sd-20;
        fc3_weights[0][11] = 16'sd-22;
        fc3_weights[0][12] = 16'sd20;
        fc3_weights[0][13] = 16'sd-43;
        fc3_weights[0][14] = 16'sd-11;
        fc3_weights[0][15] = 16'sd54;
        fc3_weights[0][16] = 16'sd-8;
        fc3_weights[0][17] = 16'sd7;
        fc3_weights[0][18] = 16'sd-10;
        fc3_weights[0][19] = 16'sd11;
        fc3_weights[0][20] = 16'sd-12;
        fc3_weights[0][21] = 16'sd-24;
        fc3_weights[0][22] = 16'sd-15;
        fc3_weights[0][23] = 16'sd-21;
        fc3_weights[0][24] = 16'sd-5;
        fc3_weights[0][25] = 16'sd0;
        fc3_weights[0][26] = 16'sd-7;
        fc3_weights[0][27] = 16'sd21;
        fc3_weights[0][28] = 16'sd14;
        fc3_weights[0][29] = 16'sd-1;
        fc3_weights[0][30] = 16'sd-1;
        fc3_weights[0][31] = 16'sd-34;
        fc3_weights[0][32] = 16'sd-2;
        fc3_weights[0][33] = 16'sd18;
        fc3_weights[0][34] = 16'sd9;
        fc3_weights[0][35] = 16'sd0;
        fc3_weights[0][36] = 16'sd-2;
        fc3_weights[0][37] = 16'sd5;
        fc3_weights[0][38] = 16'sd-3;
        fc3_weights[0][39] = 16'sd-22;
        fc3_weights[0][40] = 16'sd-47;
        fc3_weights[0][41] = 16'sd-54;
        fc3_weights[0][42] = 16'sd-2;
        fc3_weights[0][43] = 16'sd29;
        fc3_weights[0][44] = 16'sd25;
        fc3_weights[0][45] = 16'sd11;
        fc3_weights[0][46] = 16'sd3;
        fc3_weights[0][47] = 16'sd13;
        fc3_weights[0][48] = 16'sd7;
        fc3_weights[0][49] = 16'sd3;
        fc3_weights[0][50] = 16'sd-4;
        fc3_weights[0][51] = 16'sd-9;
        fc3_weights[0][52] = 16'sd3;
        fc3_weights[0][53] = 16'sd35;
        fc3_weights[0][54] = 16'sd-8;
        fc3_weights[0][55] = 16'sd-6;
        fc3_weights[0][56] = 16'sd1;
        fc3_weights[0][57] = 16'sd7;
        fc3_weights[0][58] = 16'sd10;
        fc3_weights[0][59] = 16'sd-4;
        fc3_weights[0][60] = 16'sd-10;
        fc3_weights[0][61] = 16'sd-28;
        fc3_weights[0][62] = 16'sd16;
        fc3_weights[0][63] = 16'sd1;
        fc3_weights[1][0] = 16'sd-6;
        fc3_weights[1][1] = 16'sd1;
        fc3_weights[1][2] = 16'sd-3;
        fc3_weights[1][3] = 16'sd6;
        fc3_weights[1][4] = 16'sd4;
        fc3_weights[1][5] = 16'sd-5;
        fc3_weights[1][6] = 16'sd-7;
        fc3_weights[1][7] = 16'sd3;
        fc3_weights[1][8] = 16'sd-1;
        fc3_weights[1][9] = 16'sd-1;
        fc3_weights[1][10] = 16'sd-3;
        fc3_weights[1][11] = 16'sd-4;
        fc3_weights[1][12] = 16'sd-3;
        fc3_weights[1][13] = 16'sd4;
        fc3_weights[1][14] = 16'sd3;
        fc3_weights[1][15] = 16'sd6;
        fc3_weights[1][16] = 16'sd6;
        fc3_weights[1][17] = 16'sd1;
        fc3_weights[1][18] = 16'sd-7;
        fc3_weights[1][19] = 16'sd-4;
        fc3_weights[1][20] = 16'sd-2;
        fc3_weights[1][21] = 16'sd3;
        fc3_weights[1][22] = 16'sd-3;
        fc3_weights[1][23] = 16'sd-1;
        fc3_weights[1][24] = 16'sd-1;
        fc3_weights[1][25] = 16'sd0;
        fc3_weights[1][26] = 16'sd-11;
        fc3_weights[1][27] = 16'sd-13;
        fc3_weights[1][28] = 16'sd-3;
        fc3_weights[1][29] = 16'sd6;
        fc3_weights[1][30] = 16'sd-4;
        fc3_weights[1][31] = 16'sd3;
        fc3_weights[1][32] = 16'sd-5;
        fc3_weights[1][33] = 16'sd-7;
        fc3_weights[1][34] = 16'sd1;
        fc3_weights[1][35] = 16'sd-12;
        fc3_weights[1][36] = 16'sd-5;
        fc3_weights[1][37] = 16'sd2;
        fc3_weights[1][38] = 16'sd-2;
        fc3_weights[1][39] = 16'sd5;
        fc3_weights[1][40] = 16'sd6;
        fc3_weights[1][41] = 16'sd3;
        fc3_weights[1][42] = 16'sd-1;
        fc3_weights[1][43] = 16'sd-4;
        fc3_weights[1][44] = 16'sd-4;
        fc3_weights[1][45] = 16'sd-1;
        fc3_weights[1][46] = 16'sd3;
        fc3_weights[1][47] = 16'sd-7;
        fc3_weights[1][48] = 16'sd-3;
        fc3_weights[1][49] = 16'sd2;
        fc3_weights[1][50] = 16'sd-3;
        fc3_weights[1][51] = 16'sd8;
        fc3_weights[1][52] = 16'sd-4;
        fc3_weights[1][53] = 16'sd-3;
        fc3_weights[1][54] = 16'sd0;
        fc3_weights[1][55] = 16'sd-5;
        fc3_weights[1][56] = 16'sd2;
        fc3_weights[1][57] = 16'sd-2;
        fc3_weights[1][58] = 16'sd4;
        fc3_weights[1][59] = 16'sd0;
        fc3_weights[1][60] = 16'sd-3;
        fc3_weights[1][61] = 16'sd-4;
        fc3_weights[1][62] = 16'sd-1;
        fc3_weights[1][63] = 16'sd5;
        fc3_weights[2][0] = 16'sd0;
        fc3_weights[2][1] = 16'sd-13;
        fc3_weights[2][2] = 16'sd10;
        fc3_weights[2][3] = 16'sd-6;
        fc3_weights[2][4] = 16'sd17;
        fc3_weights[2][5] = 16'sd0;
        fc3_weights[2][6] = 16'sd26;
        fc3_weights[2][7] = 16'sd-19;
        fc3_weights[2][8] = 16'sd7;
        fc3_weights[2][9] = 16'sd12;
        fc3_weights[2][10] = 16'sd-18;
        fc3_weights[2][11] = 16'sd-21;
        fc3_weights[2][12] = 16'sd18;
        fc3_weights[2][13] = 16'sd-20;
        fc3_weights[2][14] = 16'sd-17;
        fc3_weights[2][15] = 16'sd73;
        fc3_weights[2][16] = 16'sd-6;
        fc3_weights[2][17] = 16'sd9;
        fc3_weights[2][18] = 16'sd-11;
        fc3_weights[2][19] = 16'sd12;
        fc3_weights[2][20] = 16'sd-9;
        fc3_weights[2][21] = 16'sd-23;
        fc3_weights[2][22] = 16'sd-13;
        fc3_weights[2][23] = 16'sd-8;
        fc3_weights[2][24] = 16'sd-4;
        fc3_weights[2][25] = 16'sd5;
        fc3_weights[2][26] = 16'sd-8;
        fc3_weights[2][27] = 16'sd11;
        fc3_weights[2][28] = 16'sd16;
        fc3_weights[2][29] = 16'sd-3;
        fc3_weights[2][30] = 16'sd1;
        fc3_weights[2][31] = 16'sd-26;
        fc3_weights[2][32] = 16'sd-8;
        fc3_weights[2][33] = 16'sd18;
        fc3_weights[2][34] = 16'sd13;
        fc3_weights[2][35] = 16'sd-1;
        fc3_weights[2][36] = 16'sd-8;
        fc3_weights[2][37] = 16'sd0;
        fc3_weights[2][38] = 16'sd-2;
        fc3_weights[2][39] = 16'sd-13;
        fc3_weights[2][40] = 16'sd-37;
        fc3_weights[2][41] = 16'sd-50;
        fc3_weights[2][42] = 16'sd-6;
        fc3_weights[2][43] = 16'sd33;
        fc3_weights[2][44] = 16'sd22;
        fc3_weights[2][45] = 16'sd12;
        fc3_weights[2][46] = 16'sd-1;
        fc3_weights[2][47] = 16'sd3;
        fc3_weights[2][48] = 16'sd8;
        fc3_weights[2][49] = 16'sd3;
        fc3_weights[2][50] = 16'sd7;
        fc3_weights[2][51] = 16'sd-5;
        fc3_weights[2][52] = 16'sd3;
        fc3_weights[2][53] = 16'sd47;
        fc3_weights[2][54] = 16'sd-11;
        fc3_weights[2][55] = 16'sd-9;
        fc3_weights[2][56] = 16'sd8;
        fc3_weights[2][57] = 16'sd2;
        fc3_weights[2][58] = 16'sd13;
        fc3_weights[2][59] = 16'sd-6;
        fc3_weights[2][60] = 16'sd8;
        fc3_weights[2][61] = 16'sd-27;
        fc3_weights[2][62] = 16'sd21;
        fc3_weights[2][63] = 16'sd-1;
        fc3_weights[3][0] = 16'sd10;
        fc3_weights[3][1] = 16'sd-4;
        fc3_weights[3][2] = 16'sd34;
        fc3_weights[3][3] = 16'sd-12;
        fc3_weights[3][4] = 16'sd16;
        fc3_weights[3][5] = 16'sd25;
        fc3_weights[3][6] = 16'sd-17;
        fc3_weights[3][7] = 16'sd0;
        fc3_weights[3][8] = 16'sd8;
        fc3_weights[3][9] = 16'sd11;
        fc3_weights[3][10] = 16'sd5;
        fc3_weights[3][11] = 16'sd8;
        fc3_weights[3][12] = 16'sd-13;
        fc3_weights[3][13] = 16'sd62;
        fc3_weights[3][14] = 16'sd-17;
        fc3_weights[3][15] = 16'sd29;
        fc3_weights[3][16] = 16'sd-5;
        fc3_weights[3][17] = 16'sd5;
        fc3_weights[3][18] = 16'sd27;
        fc3_weights[3][19] = 16'sd11;
        fc3_weights[3][20] = 16'sd2;
        fc3_weights[3][21] = 16'sd-6;
        fc3_weights[3][22] = 16'sd-6;
        fc3_weights[3][23] = 16'sd13;
        fc3_weights[3][24] = 16'sd-2;
        fc3_weights[3][25] = 16'sd6;
        fc3_weights[3][26] = 16'sd37;
        fc3_weights[3][27] = 16'sd-5;
        fc3_weights[3][28] = 16'sd7;
        fc3_weights[3][29] = 16'sd-9;
        fc3_weights[3][30] = 16'sd8;
        fc3_weights[3][31] = 16'sd12;
        fc3_weights[3][32] = 16'sd-11;
        fc3_weights[3][33] = 16'sd22;
        fc3_weights[3][34] = 16'sd-7;
        fc3_weights[3][35] = 16'sd42;
        fc3_weights[3][36] = 16'sd-9;
        fc3_weights[3][37] = 16'sd-16;
        fc3_weights[3][38] = 16'sd-6;
        fc3_weights[3][39] = 16'sd9;
        fc3_weights[3][40] = 16'sd19;
        fc3_weights[3][41] = 16'sd11;
        fc3_weights[3][42] = 16'sd-2;
        fc3_weights[3][43] = 16'sd-22;
        fc3_weights[3][44] = 16'sd23;
        fc3_weights[3][45] = 16'sd8;
        fc3_weights[3][46] = 16'sd-9;
        fc3_weights[3][47] = 16'sd-16;
        fc3_weights[3][48] = 16'sd9;
        fc3_weights[3][49] = 16'sd-8;
        fc3_weights[3][50] = 16'sd5;
        fc3_weights[3][51] = 16'sd9;
        fc3_weights[3][52] = 16'sd13;
        fc3_weights[3][53] = 16'sd17;
        fc3_weights[3][54] = 16'sd-6;
        fc3_weights[3][55] = 16'sd26;
        fc3_weights[3][56] = 16'sd12;
        fc3_weights[3][57] = 16'sd-3;
        fc3_weights[3][58] = 16'sd0;
        fc3_weights[3][59] = 16'sd-7;
        fc3_weights[3][60] = 16'sd48;
        fc3_weights[3][61] = 16'sd8;
        fc3_weights[3][62] = 16'sd7;
        fc3_weights[3][63] = 16'sd-8;
        fc3_weights[4][0] = 16'sd44;
        fc3_weights[4][1] = 16'sd37;
        fc3_weights[4][2] = 16'sd11;
        fc3_weights[4][3] = 16'sd61;
        fc3_weights[4][4] = 16'sd15;
        fc3_weights[4][5] = 16'sd22;
        fc3_weights[4][6] = 16'sd69;
        fc3_weights[4][7] = 16'sd24;
        fc3_weights[4][8] = 16'sd187;
        fc3_weights[4][9] = 16'sd103;
        fc3_weights[4][10] = 16'sd143;
        fc3_weights[4][11] = 16'sd105;
        fc3_weights[4][12] = 16'sd158;
        fc3_weights[4][13] = 16'sd34;
        fc3_weights[4][14] = 16'sd143;
        fc3_weights[4][15] = 16'sd46;
        fc3_weights[4][16] = 16'sd159;
        fc3_weights[4][17] = 16'sd128;
        fc3_weights[4][18] = 16'sd58;
        fc3_weights[4][19] = 16'sd44;
        fc3_weights[4][20] = 16'sd77;
        fc3_weights[4][21] = 16'sd50;
        fc3_weights[4][22] = 16'sd150;
        fc3_weights[4][23] = 16'sd53;
        fc3_weights[4][24] = 16'sd170;
        fc3_weights[4][25] = 16'sd64;
        fc3_weights[4][26] = 16'sd28;
        fc3_weights[4][27] = 16'sd59;
        fc3_weights[4][28] = 16'sd79;
        fc3_weights[4][29] = 16'sd45;
        fc3_weights[4][30] = 16'sd74;
        fc3_weights[4][31] = 16'sd13;
        fc3_weights[4][32] = 16'sd127;
        fc3_weights[4][33] = 16'sd80;
        fc3_weights[4][34] = 16'sd126;
        fc3_weights[4][35] = 16'sd11;
        fc3_weights[4][36] = 16'sd70;
        fc3_weights[4][37] = 16'sd134;
        fc3_weights[4][38] = 16'sd56;
        fc3_weights[4][39] = 16'sd84;
        fc3_weights[4][40] = 16'sd50;
        fc3_weights[4][41] = 16'sd47;
        fc3_weights[4][42] = 16'sd153;
        fc3_weights[4][43] = 16'sd132;
        fc3_weights[4][44] = 16'sd37;
        fc3_weights[4][45] = 16'sd116;
        fc3_weights[4][46] = 16'sd170;
        fc3_weights[4][47] = 16'sd117;
        fc3_weights[4][48] = 16'sd145;
        fc3_weights[4][49] = 16'sd154;
        fc3_weights[4][50] = 16'sd64;
        fc3_weights[4][51] = 16'sd106;
        fc3_weights[4][52] = 16'sd38;
        fc3_weights[4][53] = 16'sd170;
        fc3_weights[4][54] = 16'sd150;
        fc3_weights[4][55] = 16'sd85;
        fc3_weights[4][56] = 16'sd12;
        fc3_weights[4][57] = 16'sd90;
        fc3_weights[4][58] = 16'sd112;
        fc3_weights[4][59] = 16'sd145;
        fc3_weights[4][60] = 16'sd6;
        fc3_weights[4][61] = 16'sd4;
        fc3_weights[4][62] = 16'sd86;
        fc3_weights[4][63] = 16'sd24;
        fc3_weights[5][0] = 16'sd-12;
        fc3_weights[5][1] = 16'sd4;
        fc3_weights[5][2] = 16'sd-2;
        fc3_weights[5][3] = 16'sd29;
        fc3_weights[5][4] = 16'sd36;
        fc3_weights[5][5] = 16'sd-33;
        fc3_weights[5][6] = 16'sd-8;
        fc3_weights[5][7] = 16'sd7;
        fc3_weights[5][8] = 16'sd-2;
        fc3_weights[5][9] = 16'sd8;
        fc3_weights[5][10] = 16'sd2;
        fc3_weights[5][11] = 16'sd-14;
        fc3_weights[5][12] = 16'sd-6;
        fc3_weights[5][13] = 16'sd-23;
        fc3_weights[5][14] = 16'sd5;
        fc3_weights[5][15] = 16'sd25;
        fc3_weights[5][16] = 16'sd14;
        fc3_weights[5][17] = 16'sd-8;
        fc3_weights[5][18] = 16'sd-26;
        fc3_weights[5][19] = 16'sd-10;
        fc3_weights[5][20] = 16'sd16;
        fc3_weights[5][21] = 16'sd-50;
        fc3_weights[5][22] = 16'sd0;
        fc3_weights[5][23] = 16'sd8;
        fc3_weights[5][24] = 16'sd-19;
        fc3_weights[5][25] = 16'sd6;
        fc3_weights[5][26] = 16'sd-49;
        fc3_weights[5][27] = 16'sd-101;
        fc3_weights[5][28] = 16'sd-11;
        fc3_weights[5][29] = 16'sd-2;
        fc3_weights[5][30] = 16'sd-9;
        fc3_weights[5][31] = 16'sd33;
        fc3_weights[5][32] = 16'sd2;
        fc3_weights[5][33] = 16'sd-62;
        fc3_weights[5][34] = 16'sd13;
        fc3_weights[5][35] = 16'sd-90;
        fc3_weights[5][36] = 16'sd15;
        fc3_weights[5][37] = 16'sd10;
        fc3_weights[5][38] = 16'sd49;
        fc3_weights[5][39] = 16'sd-6;
        fc3_weights[5][40] = 16'sd-25;
        fc3_weights[5][41] = 16'sd-42;
        fc3_weights[5][42] = 16'sd-60;
        fc3_weights[5][43] = 16'sd-49;
        fc3_weights[5][44] = 16'sd3;
        fc3_weights[5][45] = 16'sd22;
        fc3_weights[5][46] = 16'sd-1;
        fc3_weights[5][47] = 16'sd1;
        fc3_weights[5][48] = 16'sd1;
        fc3_weights[5][49] = 16'sd7;
        fc3_weights[5][50] = 16'sd-11;
        fc3_weights[5][51] = 16'sd-8;
        fc3_weights[5][52] = 16'sd-6;
        fc3_weights[5][53] = 16'sd-6;
        fc3_weights[5][54] = 16'sd-14;
        fc3_weights[5][55] = 16'sd-64;
        fc3_weights[5][56] = 16'sd-1;
        fc3_weights[5][57] = 16'sd4;
        fc3_weights[5][58] = 16'sd16;
        fc3_weights[5][59] = 16'sd17;
        fc3_weights[5][60] = 16'sd25;
        fc3_weights[5][61] = 16'sd-92;
        fc3_weights[5][62] = 16'sd22;
        fc3_weights[5][63] = 16'sd6;
        fc3_weights[6][0] = 16'sd-15;
        fc3_weights[6][1] = 16'sd2;
        fc3_weights[6][2] = 16'sd-13;
        fc3_weights[6][3] = 16'sd-8;
        fc3_weights[6][4] = 16'sd-4;
        fc3_weights[6][5] = 16'sd-17;
        fc3_weights[6][6] = 16'sd-6;
        fc3_weights[6][7] = 16'sd5;
        fc3_weights[6][8] = 16'sd3;
        fc3_weights[6][9] = 16'sd0;
        fc3_weights[6][10] = 16'sd2;
        fc3_weights[6][11] = 16'sd4;
        fc3_weights[6][12] = 16'sd3;
        fc3_weights[6][13] = 16'sd-1;
        fc3_weights[6][14] = 16'sd5;
        fc3_weights[6][15] = 16'sd-1;
        fc3_weights[6][16] = 16'sd0;
        fc3_weights[6][17] = 16'sd5;
        fc3_weights[6][18] = 16'sd-10;
        fc3_weights[6][19] = 16'sd-18;
        fc3_weights[6][20] = 16'sd-8;
        fc3_weights[6][21] = 16'sd-7;
        fc3_weights[6][22] = 16'sd1;
        fc3_weights[6][23] = 16'sd-4;
        fc3_weights[6][24] = 16'sd2;
        fc3_weights[6][25] = 16'sd-1;
        fc3_weights[6][26] = 16'sd-21;
        fc3_weights[6][27] = 16'sd0;
        fc3_weights[6][28] = 16'sd-1;
        fc3_weights[6][29] = 16'sd0;
        fc3_weights[6][30] = 16'sd0;
        fc3_weights[6][31] = 16'sd4;
        fc3_weights[6][32] = 16'sd2;
        fc3_weights[6][33] = 16'sd-25;
        fc3_weights[6][34] = 16'sd5;
        fc3_weights[6][35] = 16'sd-24;
        fc3_weights[6][36] = 16'sd-3;
        fc3_weights[6][37] = 16'sd4;
        fc3_weights[6][38] = 16'sd15;
        fc3_weights[6][39] = 16'sd3;
        fc3_weights[6][40] = 16'sd0;
        fc3_weights[6][41] = 16'sd-9;
        fc3_weights[6][42] = 16'sd-3;
        fc3_weights[6][43] = 16'sd4;
        fc3_weights[6][44] = 16'sd6;
        fc3_weights[6][45] = 16'sd3;
        fc3_weights[6][46] = 16'sd1;
        fc3_weights[6][47] = 16'sd-2;
        fc3_weights[6][48] = 16'sd3;
        fc3_weights[6][49] = 16'sd5;
        fc3_weights[6][50] = 16'sd-1;
        fc3_weights[6][51] = 16'sd2;
        fc3_weights[6][52] = 16'sd2;
        fc3_weights[6][53] = 16'sd-4;
        fc3_weights[6][54] = 16'sd4;
        fc3_weights[6][55] = 16'sd-45;
        fc3_weights[6][56] = 16'sd-5;
        fc3_weights[6][57] = 16'sd0;
        fc3_weights[6][58] = 16'sd-1;
        fc3_weights[6][59] = 16'sd10;
        fc3_weights[6][60] = 16'sd1;
        fc3_weights[6][61] = 16'sd15;
        fc3_weights[6][62] = 16'sd2;
        fc3_weights[6][63] = 16'sd6;
        fc3_weights[7][0] = 16'sd-6;
        fc3_weights[7][1] = 16'sd1;
        fc3_weights[7][2] = 16'sd-5;
        fc3_weights[7][3] = 16'sd22;
        fc3_weights[7][4] = 16'sd32;
        fc3_weights[7][5] = 16'sd-35;
        fc3_weights[7][6] = 16'sd-6;
        fc3_weights[7][7] = 16'sd1;
        fc3_weights[7][8] = 16'sd1;
        fc3_weights[7][9] = 16'sd4;
        fc3_weights[7][10] = 16'sd2;
        fc3_weights[7][11] = 16'sd-13;
        fc3_weights[7][12] = 16'sd-10;
        fc3_weights[7][13] = 16'sd-17;
        fc3_weights[7][14] = 16'sd0;
        fc3_weights[7][15] = 16'sd39;
        fc3_weights[7][16] = 16'sd11;
        fc3_weights[7][17] = 16'sd-8;
        fc3_weights[7][18] = 16'sd-21;
        fc3_weights[7][19] = 16'sd-12;
        fc3_weights[7][20] = 16'sd11;
        fc3_weights[7][21] = 16'sd-27;
        fc3_weights[7][22] = 16'sd1;
        fc3_weights[7][23] = 16'sd11;
        fc3_weights[7][24] = 16'sd-17;
        fc3_weights[7][25] = 16'sd5;
        fc3_weights[7][26] = 16'sd-47;
        fc3_weights[7][27] = 16'sd-77;
        fc3_weights[7][28] = 16'sd-10;
        fc3_weights[7][29] = 16'sd-9;
        fc3_weights[7][30] = 16'sd-5;
        fc3_weights[7][31] = 16'sd32;
        fc3_weights[7][32] = 16'sd-4;
        fc3_weights[7][33] = 16'sd-51;
        fc3_weights[7][34] = 16'sd16;
        fc3_weights[7][35] = 16'sd-69;
        fc3_weights[7][36] = 16'sd9;
        fc3_weights[7][37] = 16'sd7;
        fc3_weights[7][38] = 16'sd48;
        fc3_weights[7][39] = 16'sd-5;
        fc3_weights[7][40] = 16'sd-13;
        fc3_weights[7][41] = 16'sd-32;
        fc3_weights[7][42] = 16'sd-57;
        fc3_weights[7][43] = 16'sd-38;
        fc3_weights[7][44] = 16'sd-10;
        fc3_weights[7][45] = 16'sd20;
        fc3_weights[7][46] = 16'sd0;
        fc3_weights[7][47] = 16'sd1;
        fc3_weights[7][48] = 16'sd1;
        fc3_weights[7][49] = 16'sd7;
        fc3_weights[7][50] = 16'sd-6;
        fc3_weights[7][51] = 16'sd-13;
        fc3_weights[7][52] = 16'sd1;
        fc3_weights[7][53] = 16'sd1;
        fc3_weights[7][54] = 16'sd-12;
        fc3_weights[7][55] = 16'sd-50;
        fc3_weights[7][56] = 16'sd1;
        fc3_weights[7][57] = 16'sd3;
        fc3_weights[7][58] = 16'sd18;
        fc3_weights[7][59] = 16'sd9;
        fc3_weights[7][60] = 16'sd26;
        fc3_weights[7][61] = 16'sd-58;
        fc3_weights[7][62] = 16'sd23;
        fc3_weights[7][63] = 16'sd5;
        fc3_weights[8][0] = 16'sd30;
        fc3_weights[8][1] = 16'sd-4;
        fc3_weights[8][2] = 16'sd-12;
        fc3_weights[8][3] = 16'sd-1;
        fc3_weights[8][4] = 16'sd24;
        fc3_weights[8][5] = 16'sd28;
        fc3_weights[8][6] = 16'sd-2;
        fc3_weights[8][7] = 16'sd-10;
        fc3_weights[8][8] = 16'sd6;
        fc3_weights[8][9] = 16'sd-4;
        fc3_weights[8][10] = 16'sd1;
        fc3_weights[8][11] = 16'sd6;
        fc3_weights[8][12] = 16'sd-8;
        fc3_weights[8][13] = 16'sd10;
        fc3_weights[8][14] = 16'sd-10;
        fc3_weights[8][15] = 16'sd29;
        fc3_weights[8][16] = 16'sd-5;
        fc3_weights[8][17] = 16'sd-2;
        fc3_weights[8][18] = 16'sd21;
        fc3_weights[8][19] = 16'sd30;
        fc3_weights[8][20] = 16'sd-11;
        fc3_weights[8][21] = 16'sd17;
        fc3_weights[8][22] = 16'sd0;
        fc3_weights[8][23] = 16'sd0;
        fc3_weights[8][24] = 16'sd0;
        fc3_weights[8][25] = 16'sd-2;
        fc3_weights[8][26] = 16'sd66;
        fc3_weights[8][27] = 16'sd20;
        fc3_weights[8][28] = 16'sd1;
        fc3_weights[8][29] = 16'sd-19;
        fc3_weights[8][30] = 16'sd3;
        fc3_weights[8][31] = 16'sd-9;
        fc3_weights[8][32] = 16'sd-5;
        fc3_weights[8][33] = 16'sd29;
        fc3_weights[8][34] = 16'sd0;
        fc3_weights[8][35] = 16'sd69;
        fc3_weights[8][36] = 16'sd-10;
        fc3_weights[8][37] = 16'sd-13;
        fc3_weights[8][38] = 16'sd-3;
        fc3_weights[8][39] = 16'sd7;
        fc3_weights[8][40] = 16'sd13;
        fc3_weights[8][41] = 16'sd-5;
        fc3_weights[8][42] = 16'sd6;
        fc3_weights[8][43] = 16'sd10;
        fc3_weights[8][44] = 16'sd17;
        fc3_weights[8][45] = 16'sd-9;
        fc3_weights[8][46] = 16'sd5;
        fc3_weights[8][47] = 16'sd0;
        fc3_weights[8][48] = 16'sd4;
        fc3_weights[8][49] = 16'sd2;
        fc3_weights[8][50] = 16'sd3;
        fc3_weights[8][51] = 16'sd-5;
        fc3_weights[8][52] = 16'sd18;
        fc3_weights[8][53] = 16'sd2;
        fc3_weights[8][54] = 16'sd0;
        fc3_weights[8][55] = 16'sd68;
        fc3_weights[8][56] = 16'sd-4;
        fc3_weights[8][57] = 16'sd-3;
        fc3_weights[8][58] = 16'sd-7;
        fc3_weights[8][59] = 16'sd-16;
        fc3_weights[8][60] = 16'sd7;
        fc3_weights[8][61] = 16'sd66;
        fc3_weights[8][62] = 16'sd5;
        fc3_weights[8][63] = 16'sd0;
        fc3_weights[9][0] = 16'sd-90;
        fc3_weights[9][1] = 16'sd94;
        fc3_weights[9][2] = 16'sd56;
        fc3_weights[9][3] = 16'sd-79;
        fc3_weights[9][4] = 16'sd-59;
        fc3_weights[9][5] = 16'sd-23;
        fc3_weights[9][6] = 16'sd26;
        fc3_weights[9][7] = 16'sd67;
        fc3_weights[9][8] = 16'sd73;
        fc3_weights[9][9] = 16'sd-11;
        fc3_weights[9][10] = 16'sd58;
        fc3_weights[9][11] = 16'sd-28;
        fc3_weights[9][12] = 16'sd8;
        fc3_weights[9][13] = 16'sd7;
        fc3_weights[9][14] = 16'sd-12;
        fc3_weights[9][15] = 16'sd95;
        fc3_weights[9][16] = 16'sd8;
        fc3_weights[9][17] = 16'sd-42;
        fc3_weights[9][18] = 16'sd-52;
        fc3_weights[9][19] = 16'sd-64;
        fc3_weights[9][20] = 16'sd-81;
        fc3_weights[9][21] = 16'sd17;
        fc3_weights[9][22] = 16'sd102;
        fc3_weights[9][23] = 16'sd104;
        fc3_weights[9][24] = 16'sd100;
        fc3_weights[9][25] = 16'sd105;
        fc3_weights[9][26] = 16'sd-16;
        fc3_weights[9][27] = 16'sd27;
        fc3_weights[9][28] = 16'sd76;
        fc3_weights[9][29] = 16'sd0;
        fc3_weights[9][30] = 16'sd152;
        fc3_weights[9][31] = 16'sd-61;
        fc3_weights[9][32] = 16'sd135;
        fc3_weights[9][33] = 16'sd-29;
        fc3_weights[9][34] = 16'sd-17;
        fc3_weights[9][35] = 16'sd-33;
        fc3_weights[9][36] = 16'sd72;
        fc3_weights[9][37] = 16'sd-34;
        fc3_weights[9][38] = 16'sd-55;
        fc3_weights[9][39] = 16'sd141;
        fc3_weights[9][40] = 16'sd74;
        fc3_weights[9][41] = 16'sd18;
        fc3_weights[9][42] = 16'sd-42;
        fc3_weights[9][43] = 16'sd-29;
        fc3_weights[9][44] = 16'sd-49;
        fc3_weights[9][45] = 16'sd-39;
        fc3_weights[9][46] = 16'sd117;
        fc3_weights[9][47] = 16'sd103;
        fc3_weights[9][48] = 16'sd-32;
        fc3_weights[9][49] = 16'sd42;
        fc3_weights[9][50] = 16'sd87;
        fc3_weights[9][51] = 16'sd121;
        fc3_weights[9][52] = 16'sd-63;
        fc3_weights[9][53] = 16'sd-20;
        fc3_weights[9][54] = 16'sd88;
        fc3_weights[9][55] = 16'sd-66;
        fc3_weights[9][56] = 16'sd51;
        fc3_weights[9][57] = 16'sd95;
        fc3_weights[9][58] = 16'sd-74;
        fc3_weights[9][59] = 16'sd-67;
        fc3_weights[9][60] = 16'sd125;
        fc3_weights[9][61] = 16'sd-21;
        fc3_weights[9][62] = 16'sd83;
        fc3_weights[9][63] = 16'sd121;
        fc3_weights[10][0] = 16'sd-46;
        fc3_weights[10][1] = 16'sd-13;
        fc3_weights[10][2] = 16'sd-24;
        fc3_weights[10][3] = 16'sd6;
        fc3_weights[10][4] = 16'sd1;
        fc3_weights[10][5] = 16'sd-62;
        fc3_weights[10][6] = 16'sd12;
        fc3_weights[10][7] = 16'sd-3;
        fc3_weights[10][8] = 16'sd10;
        fc3_weights[10][9] = 16'sd-28;
        fc3_weights[10][10] = 16'sd-1;
        fc3_weights[10][11] = 16'sd-10;
        fc3_weights[10][12] = 16'sd10;
        fc3_weights[10][13] = 16'sd-38;
        fc3_weights[10][14] = 16'sd-6;
        fc3_weights[10][15] = 16'sd6;
        fc3_weights[10][16] = 16'sd29;
        fc3_weights[10][17] = 16'sd8;
        fc3_weights[10][18] = 16'sd-41;
        fc3_weights[10][19] = 16'sd-13;
        fc3_weights[10][20] = 16'sd7;
        fc3_weights[10][21] = 16'sd-14;
        fc3_weights[10][22] = 16'sd-11;
        fc3_weights[10][23] = 16'sd0;
        fc3_weights[10][24] = 16'sd-11;
        fc3_weights[10][25] = 16'sd8;
        fc3_weights[10][26] = 16'sd-44;
        fc3_weights[10][27] = 16'sd-42;
        fc3_weights[10][28] = 16'sd-13;
        fc3_weights[10][29] = 16'sd-10;
        fc3_weights[10][30] = 16'sd-10;
        fc3_weights[10][31] = 16'sd62;
        fc3_weights[10][32] = 16'sd-7;
        fc3_weights[10][33] = 16'sd-23;
        fc3_weights[10][34] = 16'sd5;
        fc3_weights[10][35] = 16'sd-43;
        fc3_weights[10][36] = 16'sd-13;
        fc3_weights[10][37] = 16'sd13;
        fc3_weights[10][38] = 16'sd18;
        fc3_weights[10][39] = 16'sd-16;
        fc3_weights[10][40] = 16'sd-27;
        fc3_weights[10][41] = 16'sd-5;
        fc3_weights[10][42] = 16'sd-36;
        fc3_weights[10][43] = 16'sd-5;
        fc3_weights[10][44] = 16'sd-11;
        fc3_weights[10][45] = 16'sd3;
        fc3_weights[10][46] = 16'sd3;
        fc3_weights[10][47] = 16'sd8;
        fc3_weights[10][48] = 16'sd-40;
        fc3_weights[10][49] = 16'sd-7;
        fc3_weights[10][50] = 16'sd7;
        fc3_weights[10][51] = 16'sd20;
        fc3_weights[10][52] = 16'sd-15;
        fc3_weights[10][53] = 16'sd17;
        fc3_weights[10][54] = 16'sd-5;
        fc3_weights[10][55] = 16'sd-51;
        fc3_weights[10][56] = 16'sd5;
        fc3_weights[10][57] = 16'sd-24;
        fc3_weights[10][58] = 16'sd6;
        fc3_weights[10][59] = 16'sd-22;
        fc3_weights[10][60] = 16'sd5;
        fc3_weights[10][61] = 16'sd-20;
        fc3_weights[10][62] = 16'sd14;
        fc3_weights[10][63] = 16'sd-7;
        fc3_weights[11][0] = 16'sd-8;
        fc3_weights[11][1] = 16'sd4;
        fc3_weights[11][2] = 16'sd-1;
        fc3_weights[11][3] = 16'sd3;
        fc3_weights[11][4] = 16'sd4;
        fc3_weights[11][5] = 16'sd2;
        fc3_weights[11][6] = 16'sd-8;
        fc3_weights[11][7] = 16'sd3;
        fc3_weights[11][8] = 16'sd-1;
        fc3_weights[11][9] = 16'sd7;
        fc3_weights[11][10] = 16'sd0;
        fc3_weights[11][11] = 16'sd5;
        fc3_weights[11][12] = 16'sd-2;
        fc3_weights[11][13] = 16'sd12;
        fc3_weights[11][14] = 16'sd2;
        fc3_weights[11][15] = 16'sd5;
        fc3_weights[11][16] = 16'sd-2;
        fc3_weights[11][17] = 16'sd5;
        fc3_weights[11][18] = 16'sd-10;
        fc3_weights[11][19] = 16'sd-1;
        fc3_weights[11][20] = 16'sd-13;
        fc3_weights[11][21] = 16'sd-1;
        fc3_weights[11][22] = 16'sd2;
        fc3_weights[11][23] = 16'sd-2;
        fc3_weights[11][24] = 16'sd0;
        fc3_weights[11][25] = 16'sd3;
        fc3_weights[11][26] = 16'sd-1;
        fc3_weights[11][27] = 16'sd5;
        fc3_weights[11][28] = 16'sd1;
        fc3_weights[11][29] = 16'sd-2;
        fc3_weights[11][30] = 16'sd-2;
        fc3_weights[11][31] = 16'sd-3;
        fc3_weights[11][32] = 16'sd2;
        fc3_weights[11][33] = 16'sd-7;
        fc3_weights[11][34] = 16'sd1;
        fc3_weights[11][35] = 16'sd4;
        fc3_weights[11][36] = 16'sd-1;
        fc3_weights[11][37] = 16'sd-2;
        fc3_weights[11][38] = 16'sd1;
        fc3_weights[11][39] = 16'sd2;
        fc3_weights[11][40] = 16'sd1;
        fc3_weights[11][41] = 16'sd-19;
        fc3_weights[11][42] = 16'sd-5;
        fc3_weights[11][43] = 16'sd0;
        fc3_weights[11][44] = 16'sd-3;
        fc3_weights[11][45] = 16'sd-3;
        fc3_weights[11][46] = 16'sd0;
        fc3_weights[11][47] = 16'sd-5;
        fc3_weights[11][48] = 16'sd3;
        fc3_weights[11][49] = 16'sd-2;
        fc3_weights[11][50] = 16'sd-4;
        fc3_weights[11][51] = 16'sd-6;
        fc3_weights[11][52] = 16'sd-2;
        fc3_weights[11][53] = 16'sd1;
        fc3_weights[11][54] = 16'sd0;
        fc3_weights[11][55] = 16'sd-4;
        fc3_weights[11][56] = 16'sd-2;
        fc3_weights[11][57] = 16'sd-1;
        fc3_weights[11][58] = 16'sd-2;
        fc3_weights[11][59] = 16'sd4;
        fc3_weights[11][60] = 16'sd-1;
        fc3_weights[11][61] = 16'sd2;
        fc3_weights[11][62] = 16'sd-2;
        fc3_weights[11][63] = 16'sd4;
        fc3_weights[12][0] = 16'sd-49;
        fc3_weights[12][1] = 16'sd-19;
        fc3_weights[12][2] = 16'sd-25;
        fc3_weights[12][3] = 16'sd2;
        fc3_weights[12][4] = 16'sd2;
        fc3_weights[12][5] = 16'sd-64;
        fc3_weights[12][6] = 16'sd15;
        fc3_weights[12][7] = 16'sd-3;
        fc3_weights[12][8] = 16'sd15;
        fc3_weights[12][9] = 16'sd-32;
        fc3_weights[12][10] = 16'sd-1;
        fc3_weights[12][11] = 16'sd-8;
        fc3_weights[12][12] = 16'sd17;
        fc3_weights[12][13] = 16'sd-44;
        fc3_weights[12][14] = 16'sd-8;
        fc3_weights[12][15] = 16'sd13;
        fc3_weights[12][16] = 16'sd25;
        fc3_weights[12][17] = 16'sd16;
        fc3_weights[12][18] = 16'sd-28;
        fc3_weights[12][19] = 16'sd-11;
        fc3_weights[12][20] = 16'sd3;
        fc3_weights[12][21] = 16'sd-5;
        fc3_weights[12][22] = 16'sd-12;
        fc3_weights[12][23] = 16'sd3;
        fc3_weights[12][24] = 16'sd-13;
        fc3_weights[12][25] = 16'sd8;
        fc3_weights[12][26] = 16'sd-50;
        fc3_weights[12][27] = 16'sd-32;
        fc3_weights[12][28] = 16'sd-16;
        fc3_weights[12][29] = 16'sd-16;
        fc3_weights[12][30] = 16'sd-10;
        fc3_weights[12][31] = 16'sd56;
        fc3_weights[12][32] = 16'sd-11;
        fc3_weights[12][33] = 16'sd-23;
        fc3_weights[12][34] = 16'sd2;
        fc3_weights[12][35] = 16'sd-49;
        fc3_weights[12][36] = 16'sd-14;
        fc3_weights[12][37] = 16'sd17;
        fc3_weights[12][38] = 16'sd21;
        fc3_weights[12][39] = 16'sd-14;
        fc3_weights[12][40] = 16'sd-25;
        fc3_weights[12][41] = 16'sd7;
        fc3_weights[12][42] = 16'sd-30;
        fc3_weights[12][43] = 16'sd-5;
        fc3_weights[12][44] = 16'sd-13;
        fc3_weights[12][45] = 16'sd1;
        fc3_weights[12][46] = 16'sd1;
        fc3_weights[12][47] = 16'sd6;
        fc3_weights[12][48] = 16'sd-34;
        fc3_weights[12][49] = 16'sd-9;
        fc3_weights[12][50] = 16'sd8;
        fc3_weights[12][51] = 16'sd16;
        fc3_weights[12][52] = 16'sd-23;
        fc3_weights[12][53] = 16'sd21;
        fc3_weights[12][54] = 16'sd-1;
        fc3_weights[12][55] = 16'sd-44;
        fc3_weights[12][56] = 16'sd6;
        fc3_weights[12][57] = 16'sd-20;
        fc3_weights[12][58] = 16'sd14;
        fc3_weights[12][59] = 16'sd-12;
        fc3_weights[12][60] = 16'sd8;
        fc3_weights[12][61] = 16'sd-17;
        fc3_weights[12][62] = 16'sd16;
        fc3_weights[12][63] = 16'sd-9;
        fc3_weights[13][0] = 16'sd32;
        fc3_weights[13][1] = 16'sd6;
        fc3_weights[13][2] = 16'sd0;
        fc3_weights[13][3] = 16'sd8;
        fc3_weights[13][4] = 16'sd19;
        fc3_weights[13][5] = 16'sd22;
        fc3_weights[13][6] = 16'sd-7;
        fc3_weights[13][7] = 16'sd3;
        fc3_weights[13][8] = 16'sd6;
        fc3_weights[13][9] = 16'sd12;
        fc3_weights[13][10] = 16'sd0;
        fc3_weights[13][11] = 16'sd6;
        fc3_weights[13][12] = 16'sd-7;
        fc3_weights[13][13] = 16'sd12;
        fc3_weights[13][14] = 16'sd-13;
        fc3_weights[13][15] = 16'sd25;
        fc3_weights[13][16] = 16'sd-4;
        fc3_weights[13][17] = 16'sd0;
        fc3_weights[13][18] = 16'sd28;
        fc3_weights[13][19] = 16'sd18;
        fc3_weights[13][20] = 16'sd-10;
        fc3_weights[13][21] = 16'sd10;
        fc3_weights[13][22] = 16'sd-4;
        fc3_weights[13][23] = 16'sd-1;
        fc3_weights[13][24] = 16'sd-3;
        fc3_weights[13][25] = 16'sd2;
        fc3_weights[13][26] = 16'sd52;
        fc3_weights[13][27] = 16'sd9;
        fc3_weights[13][28] = 16'sd5;
        fc3_weights[13][29] = 16'sd9;
        fc3_weights[13][30] = 16'sd-5;
        fc3_weights[13][31] = 16'sd-2;
        fc3_weights[13][32] = 16'sd0;
        fc3_weights[13][33] = 16'sd35;
        fc3_weights[13][34] = 16'sd-1;
        fc3_weights[13][35] = 16'sd30;
        fc3_weights[13][36] = 16'sd-1;
        fc3_weights[13][37] = 16'sd-13;
        fc3_weights[13][38] = 16'sd16;
        fc3_weights[13][39] = 16'sd3;
        fc3_weights[13][40] = 16'sd17;
        fc3_weights[13][41] = 16'sd-4;
        fc3_weights[13][42] = 16'sd7;
        fc3_weights[13][43] = 16'sd-5;
        fc3_weights[13][44] = 16'sd8;
        fc3_weights[13][45] = 16'sd-3;
        fc3_weights[13][46] = 16'sd5;
        fc3_weights[13][47] = 16'sd0;
        fc3_weights[13][48] = 16'sd16;
        fc3_weights[13][49] = 16'sd-6;
        fc3_weights[13][50] = 16'sd-1;
        fc3_weights[13][51] = 16'sd-4;
        fc3_weights[13][52] = 16'sd23;
        fc3_weights[13][53] = 16'sd9;
        fc3_weights[13][54] = 16'sd3;
        fc3_weights[13][55] = 16'sd17;
        fc3_weights[13][56] = 16'sd-3;
        fc3_weights[13][57] = 16'sd0;
        fc3_weights[13][58] = 16'sd-8;
        fc3_weights[13][59] = 16'sd13;
        fc3_weights[13][60] = 16'sd-5;
        fc3_weights[13][61] = 16'sd38;
        fc3_weights[13][62] = 16'sd5;
        fc3_weights[13][63] = 16'sd-4;
        fc3_weights[14][0] = 16'sd-108;
        fc3_weights[14][1] = 16'sd-84;
        fc3_weights[14][2] = 16'sd-140;
        fc3_weights[14][3] = 16'sd-82;
        fc3_weights[14][4] = 16'sd-48;
        fc3_weights[14][5] = 16'sd-14;
        fc3_weights[14][6] = 16'sd60;
        fc3_weights[14][7] = 16'sd-114;
        fc3_weights[14][8] = 16'sd-1;
        fc3_weights[14][9] = 16'sd-112;
        fc3_weights[14][10] = 16'sd79;
        fc3_weights[14][11] = 16'sd-75;
        fc3_weights[14][12] = 16'sd-63;
        fc3_weights[14][13] = 16'sd23;
        fc3_weights[14][14] = 16'sd-98;
        fc3_weights[14][15] = 16'sd4;
        fc3_weights[14][16] = 16'sd-46;
        fc3_weights[14][17] = 16'sd-60;
        fc3_weights[14][18] = 16'sd-82;
        fc3_weights[14][19] = 16'sd-42;
        fc3_weights[14][20] = 16'sd-100;
        fc3_weights[14][21] = 16'sd-91;
        fc3_weights[14][22] = 16'sd-33;
        fc3_weights[14][23] = 16'sd80;
        fc3_weights[14][24] = 16'sd-38;
        fc3_weights[14][25] = 16'sd63;
        fc3_weights[14][26] = 16'sd-76;
        fc3_weights[14][27] = 16'sd8;
        fc3_weights[14][28] = 16'sd-46;
        fc3_weights[14][29] = 16'sd-94;
        fc3_weights[14][30] = 16'sd77;
        fc3_weights[14][31] = 16'sd32;
        fc3_weights[14][32] = 16'sd18;
        fc3_weights[14][33] = 16'sd-86;
        fc3_weights[14][34] = 16'sd-92;
        fc3_weights[14][35] = 16'sd-49;
        fc3_weights[14][36] = 16'sd49;
        fc3_weights[14][37] = 16'sd-65;
        fc3_weights[14][38] = 16'sd-56;
        fc3_weights[14][39] = 16'sd-17;
        fc3_weights[14][40] = 16'sd-36;
        fc3_weights[14][41] = 16'sd-17;
        fc3_weights[14][42] = 16'sd48;
        fc3_weights[14][43] = 16'sd-4;
        fc3_weights[14][44] = 16'sd-1;
        fc3_weights[14][45] = 16'sd-63;
        fc3_weights[14][46] = 16'sd32;
        fc3_weights[14][47] = 16'sd39;
        fc3_weights[14][48] = 16'sd-118;
        fc3_weights[14][49] = 16'sd-83;
        fc3_weights[14][50] = 16'sd115;
        fc3_weights[14][51] = 16'sd55;
        fc3_weights[14][52] = 16'sd-84;
        fc3_weights[14][53] = 16'sd-39;
        fc3_weights[14][54] = 16'sd69;
        fc3_weights[14][55] = 16'sd4;
        fc3_weights[14][56] = 16'sd-105;
        fc3_weights[14][57] = 16'sd-66;
        fc3_weights[14][58] = 16'sd-31;
        fc3_weights[14][59] = 16'sd-85;
        fc3_weights[14][60] = 16'sd-16;
        fc3_weights[14][61] = 16'sd-96;
        fc3_weights[14][62] = 16'sd34;
        fc3_weights[14][63] = 16'sd63;
        // fc3 biases
        fc3_biases[0] = 16'sd-44;
        fc3_biases[1] = 16'sd-54;
        fc3_biases[2] = 16'sd18;
        fc3_biases[3] = 16'sd111;
        fc3_biases[4] = 16'sd139;
        fc3_biases[5] = 16'sd-21;
        fc3_biases[6] = 16'sd-63;
        fc3_biases[7] = 16'sd16;
        fc3_biases[8] = 16'sd24;
        fc3_biases[9] = 16'sd47;
        fc3_biases[10] = 16'sd-2;
        fc3_biases[11] = 16'sd-58;
        fc3_biases[12] = 16'sd26;
        fc3_biases[13] = 16'sd-8;
        fc3_biases[14] = 16'sd-8;
        
        
    end

endmodule
